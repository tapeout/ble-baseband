`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module ble_crc(
  input         clock,
  input         reset,
  input         io_operand_valid,
  input         io_operand_bits,
  output [23:0] io_result_bits,
  input  [23:0] io_seed,
  input         io_init
);
  reg [23:0] lfsr; // @[Serial_CRC.scala 73:19]
  reg [31:0] _RAND_0;
  wire  _T_18; // @[Serial_CRC.scala 74:20]
  wire  inv; // @[Serial_CRC.scala 74:24]
  wire [15:0] _T_22; // @[Bitwise.scala 109:18]
  wire [7:0] _T_27; // @[Bitwise.scala 103:21]
  wire [15:0] _T_28; // @[Bitwise.scala 103:31]
  wire [7:0] _T_29; // @[Bitwise.scala 103:46]
  wire [15:0] _GEN_4; // @[Bitwise.scala 103:65]
  wire [15:0] _T_30; // @[Bitwise.scala 103:65]
  wire [15:0] _T_32; // @[Bitwise.scala 103:75]
  wire [15:0] _T_33; // @[Bitwise.scala 103:39]
  wire [11:0] _T_37; // @[Bitwise.scala 103:21]
  wire [15:0] _GEN_5; // @[Bitwise.scala 103:31]
  wire [15:0] _T_38; // @[Bitwise.scala 103:31]
  wire [11:0] _T_39; // @[Bitwise.scala 103:46]
  wire [15:0] _GEN_6; // @[Bitwise.scala 103:65]
  wire [15:0] _T_40; // @[Bitwise.scala 103:65]
  wire [15:0] _T_42; // @[Bitwise.scala 103:75]
  wire [15:0] _T_43; // @[Bitwise.scala 103:39]
  wire [13:0] _T_47; // @[Bitwise.scala 103:21]
  wire [15:0] _GEN_7; // @[Bitwise.scala 103:31]
  wire [15:0] _T_48; // @[Bitwise.scala 103:31]
  wire [13:0] _T_49; // @[Bitwise.scala 103:46]
  wire [15:0] _GEN_8; // @[Bitwise.scala 103:65]
  wire [15:0] _T_50; // @[Bitwise.scala 103:65]
  wire [15:0] _T_52; // @[Bitwise.scala 103:75]
  wire [15:0] _T_53; // @[Bitwise.scala 103:39]
  wire [14:0] _T_57; // @[Bitwise.scala 103:21]
  wire [15:0] _GEN_9; // @[Bitwise.scala 103:31]
  wire [15:0] _T_58; // @[Bitwise.scala 103:31]
  wire [14:0] _T_59; // @[Bitwise.scala 103:46]
  wire [15:0] _GEN_10; // @[Bitwise.scala 103:65]
  wire [15:0] _T_60; // @[Bitwise.scala 103:65]
  wire [15:0] _T_62; // @[Bitwise.scala 103:75]
  wire [15:0] _T_63; // @[Bitwise.scala 103:39]
  wire [7:0] _T_64; // @[Bitwise.scala 109:44]
  wire [3:0] _T_69; // @[Bitwise.scala 103:21]
  wire [7:0] _T_70; // @[Bitwise.scala 103:31]
  wire [3:0] _T_71; // @[Bitwise.scala 103:46]
  wire [7:0] _GEN_11; // @[Bitwise.scala 103:65]
  wire [7:0] _T_72; // @[Bitwise.scala 103:65]
  wire [7:0] _T_74; // @[Bitwise.scala 103:75]
  wire [7:0] _T_75; // @[Bitwise.scala 103:39]
  wire [5:0] _T_79; // @[Bitwise.scala 103:21]
  wire [7:0] _GEN_12; // @[Bitwise.scala 103:31]
  wire [7:0] _T_80; // @[Bitwise.scala 103:31]
  wire [5:0] _T_81; // @[Bitwise.scala 103:46]
  wire [7:0] _GEN_13; // @[Bitwise.scala 103:65]
  wire [7:0] _T_82; // @[Bitwise.scala 103:65]
  wire [7:0] _T_84; // @[Bitwise.scala 103:75]
  wire [7:0] _T_85; // @[Bitwise.scala 103:39]
  wire [6:0] _T_89; // @[Bitwise.scala 103:21]
  wire [7:0] _GEN_14; // @[Bitwise.scala 103:31]
  wire [7:0] _T_90; // @[Bitwise.scala 103:31]
  wire [6:0] _T_91; // @[Bitwise.scala 103:46]
  wire [7:0] _GEN_15; // @[Bitwise.scala 103:65]
  wire [7:0] _T_92; // @[Bitwise.scala 103:65]
  wire [7:0] _T_94; // @[Bitwise.scala 103:75]
  wire [7:0] _T_95; // @[Bitwise.scala 103:39]
  wire [23:0] _T_96; // @[Cat.scala 30:58]
  wire  _T_101; // @[Serial_CRC.scala 95:28]
  wire  _T_102; // @[Serial_CRC.scala 95:32]
  wire  _T_103; // @[Serial_CRC.scala 95:42]
  wire  _T_104; // @[Serial_CRC.scala 95:51]
  wire  _T_105; // @[Serial_CRC.scala 95:55]
  wire  _T_106; // @[Serial_CRC.scala 95:64]
  wire  _T_107; // @[Serial_CRC.scala 95:68]
  wire  _T_108; // @[Serial_CRC.scala 95:77]
  wire  _T_109; // @[Serial_CRC.scala 95:86]
  wire  _T_110; // @[Serial_CRC.scala 95:90]
  wire  _T_111; // @[Serial_CRC.scala 95:100]
  wire  _T_112; // @[Serial_CRC.scala 96:13]
  wire  _T_113; // @[Serial_CRC.scala 96:22]
  wire  _T_114; // @[Serial_CRC.scala 96:26]
  wire  _T_115; // @[Serial_CRC.scala 96:35]
  wire  _T_116; // @[Serial_CRC.scala 96:39]
  wire  _T_117; // @[Serial_CRC.scala 96:48]
  wire  _T_118; // @[Serial_CRC.scala 96:57]
  wire  _T_119; // @[Serial_CRC.scala 96:66]
  wire  _T_120; // @[Serial_CRC.scala 96:75]
  wire  _T_121; // @[Serial_CRC.scala 96:84]
  wire  _T_122; // @[Serial_CRC.scala 96:92]
  wire  _T_123; // @[Serial_CRC.scala 97:13]
  wire  _T_124; // @[Serial_CRC.scala 97:22]
  wire  _T_125; // @[Serial_CRC.scala 97:30]
  wire  _T_126; // @[Serial_CRC.scala 97:38]
  wire  _T_127; // @[Serial_CRC.scala 97:46]
  wire  _T_128; // @[Serial_CRC.scala 97:54]
  wire  _T_129; // @[Serial_CRC.scala 97:62]
  wire [1:0] _T_130; // @[Cat.scala 30:58]
  wire [2:0] _T_131; // @[Cat.scala 30:58]
  wire [1:0] _T_132; // @[Cat.scala 30:58]
  wire [2:0] _T_133; // @[Cat.scala 30:58]
  wire [5:0] _T_134; // @[Cat.scala 30:58]
  wire [1:0] _T_135; // @[Cat.scala 30:58]
  wire [2:0] _T_136; // @[Cat.scala 30:58]
  wire [1:0] _T_137; // @[Cat.scala 30:58]
  wire [2:0] _T_138; // @[Cat.scala 30:58]
  wire [5:0] _T_139; // @[Cat.scala 30:58]
  wire [11:0] _T_140; // @[Cat.scala 30:58]
  wire [1:0] _T_141; // @[Cat.scala 30:58]
  wire [2:0] _T_142; // @[Cat.scala 30:58]
  wire [1:0] _T_143; // @[Cat.scala 30:58]
  wire [2:0] _T_144; // @[Cat.scala 30:58]
  wire [5:0] _T_145; // @[Cat.scala 30:58]
  wire [1:0] _T_146; // @[Cat.scala 30:58]
  wire [2:0] _T_147; // @[Cat.scala 30:58]
  wire [1:0] _T_148; // @[Cat.scala 30:58]
  wire [2:0] _T_149; // @[Cat.scala 30:58]
  wire [5:0] _T_150; // @[Cat.scala 30:58]
  wire [11:0] _T_151; // @[Cat.scala 30:58]
  wire [23:0] _T_152; // @[Cat.scala 30:58]
  wire [23:0] _GEN_0; // @[Serial_CRC.scala 91:47]
  wire [23:0] _GEN_2; // @[Serial_CRC.scala 85:31]
  assign _T_18 = lfsr[0]; // @[Serial_CRC.scala 74:20]
  assign inv = _T_18 ^ io_operand_bits; // @[Serial_CRC.scala 74:24]
  assign _T_22 = io_seed[15:0]; // @[Bitwise.scala 109:18]
  assign _T_27 = _T_22[15:8]; // @[Bitwise.scala 103:21]
  assign _T_28 = {{8'd0}, _T_27}; // @[Bitwise.scala 103:31]
  assign _T_29 = _T_22[7:0]; // @[Bitwise.scala 103:46]
  assign _GEN_4 = {{8'd0}, _T_29}; // @[Bitwise.scala 103:65]
  assign _T_30 = _GEN_4 << 8; // @[Bitwise.scala 103:65]
  assign _T_32 = _T_30 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _T_33 = _T_28 | _T_32; // @[Bitwise.scala 103:39]
  assign _T_37 = _T_33[15:4]; // @[Bitwise.scala 103:21]
  assign _GEN_5 = {{4'd0}, _T_37}; // @[Bitwise.scala 103:31]
  assign _T_38 = _GEN_5 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _T_39 = _T_33[11:0]; // @[Bitwise.scala 103:46]
  assign _GEN_6 = {{4'd0}, _T_39}; // @[Bitwise.scala 103:65]
  assign _T_40 = _GEN_6 << 4; // @[Bitwise.scala 103:65]
  assign _T_42 = _T_40 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _T_43 = _T_38 | _T_42; // @[Bitwise.scala 103:39]
  assign _T_47 = _T_43[15:2]; // @[Bitwise.scala 103:21]
  assign _GEN_7 = {{2'd0}, _T_47}; // @[Bitwise.scala 103:31]
  assign _T_48 = _GEN_7 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _T_49 = _T_43[13:0]; // @[Bitwise.scala 103:46]
  assign _GEN_8 = {{2'd0}, _T_49}; // @[Bitwise.scala 103:65]
  assign _T_50 = _GEN_8 << 2; // @[Bitwise.scala 103:65]
  assign _T_52 = _T_50 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _T_53 = _T_48 | _T_52; // @[Bitwise.scala 103:39]
  assign _T_57 = _T_53[15:1]; // @[Bitwise.scala 103:21]
  assign _GEN_9 = {{1'd0}, _T_57}; // @[Bitwise.scala 103:31]
  assign _T_58 = _GEN_9 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _T_59 = _T_53[14:0]; // @[Bitwise.scala 103:46]
  assign _GEN_10 = {{1'd0}, _T_59}; // @[Bitwise.scala 103:65]
  assign _T_60 = _GEN_10 << 1; // @[Bitwise.scala 103:65]
  assign _T_62 = _T_60 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign _T_63 = _T_58 | _T_62; // @[Bitwise.scala 103:39]
  assign _T_64 = io_seed[23:16]; // @[Bitwise.scala 109:44]
  assign _T_69 = _T_64[7:4]; // @[Bitwise.scala 103:21]
  assign _T_70 = {{4'd0}, _T_69}; // @[Bitwise.scala 103:31]
  assign _T_71 = _T_64[3:0]; // @[Bitwise.scala 103:46]
  assign _GEN_11 = {{4'd0}, _T_71}; // @[Bitwise.scala 103:65]
  assign _T_72 = _GEN_11 << 4; // @[Bitwise.scala 103:65]
  assign _T_74 = _T_72 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _T_75 = _T_70 | _T_74; // @[Bitwise.scala 103:39]
  assign _T_79 = _T_75[7:2]; // @[Bitwise.scala 103:21]
  assign _GEN_12 = {{2'd0}, _T_79}; // @[Bitwise.scala 103:31]
  assign _T_80 = _GEN_12 & 8'h33; // @[Bitwise.scala 103:31]
  assign _T_81 = _T_75[5:0]; // @[Bitwise.scala 103:46]
  assign _GEN_13 = {{2'd0}, _T_81}; // @[Bitwise.scala 103:65]
  assign _T_82 = _GEN_13 << 2; // @[Bitwise.scala 103:65]
  assign _T_84 = _T_82 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _T_85 = _T_80 | _T_84; // @[Bitwise.scala 103:39]
  assign _T_89 = _T_85[7:1]; // @[Bitwise.scala 103:21]
  assign _GEN_14 = {{1'd0}, _T_89}; // @[Bitwise.scala 103:31]
  assign _T_90 = _GEN_14 & 8'h55; // @[Bitwise.scala 103:31]
  assign _T_91 = _T_85[6:0]; // @[Bitwise.scala 103:46]
  assign _GEN_15 = {{1'd0}, _T_91}; // @[Bitwise.scala 103:65]
  assign _T_92 = _GEN_15 << 1; // @[Bitwise.scala 103:65]
  assign _T_94 = _T_92 & 8'haa; // @[Bitwise.scala 103:75]
  assign _T_95 = _T_90 | _T_94; // @[Bitwise.scala 103:39]
  assign _T_96 = {_T_63,_T_95}; // @[Cat.scala 30:58]
  assign _T_101 = lfsr[23]; // @[Serial_CRC.scala 95:28]
  assign _T_102 = _T_101 ^ inv; // @[Serial_CRC.scala 95:32]
  assign _T_103 = lfsr[22]; // @[Serial_CRC.scala 95:42]
  assign _T_104 = lfsr[21]; // @[Serial_CRC.scala 95:51]
  assign _T_105 = _T_104 ^ inv; // @[Serial_CRC.scala 95:55]
  assign _T_106 = lfsr[20]; // @[Serial_CRC.scala 95:64]
  assign _T_107 = _T_106 ^ inv; // @[Serial_CRC.scala 95:68]
  assign _T_108 = lfsr[19]; // @[Serial_CRC.scala 95:77]
  assign _T_109 = lfsr[18]; // @[Serial_CRC.scala 95:86]
  assign _T_110 = _T_109 ^ inv; // @[Serial_CRC.scala 95:90]
  assign _T_111 = lfsr[17]; // @[Serial_CRC.scala 95:100]
  assign _T_112 = lfsr[16]; // @[Serial_CRC.scala 96:13]
  assign _T_113 = lfsr[15]; // @[Serial_CRC.scala 96:22]
  assign _T_114 = _T_113 ^ inv; // @[Serial_CRC.scala 96:26]
  assign _T_115 = lfsr[14]; // @[Serial_CRC.scala 96:35]
  assign _T_116 = _T_115 ^ inv; // @[Serial_CRC.scala 96:39]
  assign _T_117 = lfsr[13]; // @[Serial_CRC.scala 96:48]
  assign _T_118 = lfsr[12]; // @[Serial_CRC.scala 96:57]
  assign _T_119 = lfsr[11]; // @[Serial_CRC.scala 96:66]
  assign _T_120 = lfsr[10]; // @[Serial_CRC.scala 96:75]
  assign _T_121 = lfsr[9]; // @[Serial_CRC.scala 96:84]
  assign _T_122 = lfsr[8]; // @[Serial_CRC.scala 96:92]
  assign _T_123 = lfsr[7]; // @[Serial_CRC.scala 97:13]
  assign _T_124 = lfsr[6]; // @[Serial_CRC.scala 97:22]
  assign _T_125 = lfsr[5]; // @[Serial_CRC.scala 97:30]
  assign _T_126 = lfsr[4]; // @[Serial_CRC.scala 97:38]
  assign _T_127 = lfsr[3]; // @[Serial_CRC.scala 97:46]
  assign _T_128 = lfsr[2]; // @[Serial_CRC.scala 97:54]
  assign _T_129 = lfsr[1]; // @[Serial_CRC.scala 97:62]
  assign _T_130 = {_T_127,_T_128}; // @[Cat.scala 30:58]
  assign _T_131 = {_T_130,_T_129}; // @[Cat.scala 30:58]
  assign _T_132 = {_T_124,_T_125}; // @[Cat.scala 30:58]
  assign _T_133 = {_T_132,_T_126}; // @[Cat.scala 30:58]
  assign _T_134 = {_T_133,_T_131}; // @[Cat.scala 30:58]
  assign _T_135 = {_T_121,_T_122}; // @[Cat.scala 30:58]
  assign _T_136 = {_T_135,_T_123}; // @[Cat.scala 30:58]
  assign _T_137 = {_T_118,_T_119}; // @[Cat.scala 30:58]
  assign _T_138 = {_T_137,_T_120}; // @[Cat.scala 30:58]
  assign _T_139 = {_T_138,_T_136}; // @[Cat.scala 30:58]
  assign _T_140 = {_T_139,_T_134}; // @[Cat.scala 30:58]
  assign _T_141 = {_T_114,_T_116}; // @[Cat.scala 30:58]
  assign _T_142 = {_T_141,_T_117}; // @[Cat.scala 30:58]
  assign _T_143 = {_T_110,_T_111}; // @[Cat.scala 30:58]
  assign _T_144 = {_T_143,_T_112}; // @[Cat.scala 30:58]
  assign _T_145 = {_T_144,_T_142}; // @[Cat.scala 30:58]
  assign _T_146 = {_T_105,_T_107}; // @[Cat.scala 30:58]
  assign _T_147 = {_T_146,_T_108}; // @[Cat.scala 30:58]
  assign _T_148 = {inv,_T_102}; // @[Cat.scala 30:58]
  assign _T_149 = {_T_148,_T_103}; // @[Cat.scala 30:58]
  assign _T_150 = {_T_149,_T_147}; // @[Cat.scala 30:58]
  assign _T_151 = {_T_150,_T_145}; // @[Cat.scala 30:58]
  assign _T_152 = {_T_151,_T_140}; // @[Cat.scala 30:58]
  assign _GEN_0 = io_operand_valid ? _T_152 : lfsr; // @[Serial_CRC.scala 91:47]
  assign _GEN_2 = io_init ? _T_96 : _GEN_0; // @[Serial_CRC.scala 85:31]
  assign io_result_bits = lfsr;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  lfsr = _RAND_0[23:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      lfsr <= 24'h0;
    end else begin
      if (io_init) begin
        lfsr <= _T_96;
      end else begin
        if (io_operand_valid) begin
          lfsr <= _T_152;
        end
      end
    end
  end
endmodule
module ble_whitening(
  input        clock,
  input        reset,
  input        io_operand_valid,
  input        io_operand_bits,
  output       io_result_bits,
  input  [6:0] io_seed,
  input        io_init
);
  reg [6:0] whitening_lfsr; // @[whitening.scala 47:29]
  reg [31:0] _RAND_0;
  wire  inv; // @[whitening.scala 48:39]
  wire  _T_29; // @[whitening.scala 68:50]
  wire  _T_30; // @[whitening.scala 68:69]
  wire  _T_31; // @[whitening.scala 68:87]
  wire  _T_32; // @[whitening.scala 68:105]
  wire  _T_33; // @[whitening.scala 68:108]
  wire  _T_34; // @[whitening.scala 68:127]
  wire  _T_35; // @[whitening.scala 68:145]
  wire [1:0] _T_36; // @[Cat.scala 30:58]
  wire [2:0] _T_37; // @[Cat.scala 30:58]
  wire [1:0] _T_38; // @[Cat.scala 30:58]
  wire [1:0] _T_39; // @[Cat.scala 30:58]
  wire [3:0] _T_40; // @[Cat.scala 30:58]
  wire [6:0] _T_41; // @[Cat.scala 30:58]
  wire  _T_42; // @[whitening.scala 72:27]
  wire [6:0] _GEN_0; // @[whitening.scala 67:47]
  wire  _GEN_1; // @[whitening.scala 67:47]
  wire [6:0] _GEN_3; // @[whitening.scala 59:31]
  wire  output_bit; // @[whitening.scala 59:31]
  assign inv = whitening_lfsr[0]; // @[whitening.scala 48:39]
  assign _T_29 = whitening_lfsr[6]; // @[whitening.scala 68:50]
  assign _T_30 = whitening_lfsr[5]; // @[whitening.scala 68:69]
  assign _T_31 = whitening_lfsr[4]; // @[whitening.scala 68:87]
  assign _T_32 = whitening_lfsr[3]; // @[whitening.scala 68:105]
  assign _T_33 = _T_32 ^ inv; // @[whitening.scala 68:108]
  assign _T_34 = whitening_lfsr[2]; // @[whitening.scala 68:127]
  assign _T_35 = whitening_lfsr[1]; // @[whitening.scala 68:145]
  assign _T_36 = {_T_33,_T_34}; // @[Cat.scala 30:58]
  assign _T_37 = {_T_36,_T_35}; // @[Cat.scala 30:58]
  assign _T_38 = {_T_30,_T_31}; // @[Cat.scala 30:58]
  assign _T_39 = {inv,_T_29}; // @[Cat.scala 30:58]
  assign _T_40 = {_T_39,_T_38}; // @[Cat.scala 30:58]
  assign _T_41 = {_T_40,_T_37}; // @[Cat.scala 30:58]
  assign _T_42 = inv ^ io_operand_bits; // @[whitening.scala 72:27]
  assign _GEN_0 = io_operand_valid ? _T_41 : whitening_lfsr; // @[whitening.scala 67:47]
  assign _GEN_1 = io_operand_valid ? _T_42 : 1'h0; // @[whitening.scala 67:47]
  assign _GEN_3 = io_init ? io_seed : _GEN_0; // @[whitening.scala 59:31]
  assign output_bit = io_init ? 1'h0 : _GEN_1; // @[whitening.scala 59:31]
  assign io_result_bits = output_bit;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  whitening_lfsr = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      whitening_lfsr <= 7'h0;
    end else begin
      if (io_init) begin
        whitening_lfsr <= io_seed;
      end else begin
        if (io_operand_valid) begin
          whitening_lfsr <= _T_41;
        end
      end
    end
  end
endmodule
module ble_packetdisassembler(
  input         clock,
  input         reset,
  input         io_DMA_Switch_i,
  input  [31:0] io_REG_AA_i,
  input  [23:0] io_REG_CRC_Seed_i,
  input  [6:0]  io_REG_DeWhite_Seed_i,
  input         io_DMA_Data_o_ready,
  output        io_DMA_Data_o_valid,
  output [7:0]  io_DMA_Data_o_bits,
  input         io_DMA_Length_o_ready,
  output        io_DMA_Length_o_valid,
  output [7:0]  io_DMA_Length_o_bits,
  input         io_DMA_Flag_AA_o_ready,
  output        io_DMA_Flag_AA_o_valid,
  output        io_DMA_Flag_AA_o_bits,
  input         io_DMA_Flag_CRC_o_ready,
  output        io_DMA_Flag_CRC_o_valid,
  output        io_DMA_Flag_CRC_o_bits,
  output        io_AFIFO_Data_i_ready,
  input         io_AFIFO_Data_i_valid,
  input         io_AFIFO_Data_i_bits
);
  reg [2:0] state_r; // @[disassembler.scala 65:24]
  reg [31:0] _RAND_0;
  reg [7:0] counter_r; // @[disassembler.scala 68:26]
  reg [31:0] _RAND_1;
  reg [2:0] counter_byte_r; // @[disassembler.scala 71:31]
  reg [31:0] _RAND_2;
  reg [7:0] PDU_Length_r; // @[disassembler.scala 74:29]
  reg [31:0] _RAND_3;
  reg  PDU_Length_Valid_r; // @[disassembler.scala 75:35]
  reg [31:0] _RAND_4;
  reg  Flag_AA_r; // @[disassembler.scala 76:26]
  reg [31:0] _RAND_5;
  reg  Flag_AA_Valid_r; // @[disassembler.scala 77:32]
  reg [31:0] _RAND_6;
  reg  Flag_CRC_r; // @[disassembler.scala 78:27]
  reg [31:0] _RAND_7;
  reg  Flag_CRC_Valid_r; // @[disassembler.scala 79:33]
  reg [31:0] _RAND_8;
  reg  DMA_Data_Valid_r; // @[disassembler.scala 87:33]
  reg [31:0] _RAND_9;
  reg  AFIFO_Ready_r; // @[disassembler.scala 91:30]
  reg [31:0] _RAND_10;
  reg [7:0] data_r; // @[disassembler.scala 97:23]
  reg [31:0] _RAND_11;
  wire  CRC_inst_clock; // @[disassembler.scala 425:24]
  wire  CRC_inst_reset; // @[disassembler.scala 425:24]
  wire  CRC_inst_io_operand_valid; // @[disassembler.scala 425:24]
  wire  CRC_inst_io_operand_bits; // @[disassembler.scala 425:24]
  wire [23:0] CRC_inst_io_result_bits; // @[disassembler.scala 425:24]
  wire [23:0] CRC_inst_io_seed; // @[disassembler.scala 425:24]
  wire  CRC_inst_io_init; // @[disassembler.scala 425:24]
  wire  WHITE_inst_clock; // @[disassembler.scala 435:26]
  wire  WHITE_inst_reset; // @[disassembler.scala 435:26]
  wire  WHITE_inst_io_operand_valid; // @[disassembler.scala 435:26]
  wire  WHITE_inst_io_operand_bits; // @[disassembler.scala 435:26]
  wire  WHITE_inst_io_result_bits; // @[disassembler.scala 435:26]
  wire [6:0] WHITE_inst_io_seed; // @[disassembler.scala 435:26]
  wire  WHITE_inst_io_init; // @[disassembler.scala 435:26]
  wire  DMA_Data_Fire_w; // @[disassembler.scala 115:42]
  wire  AFIFO_Fire_w; // @[disassembler.scala 116:41]
  wire  _T_102; // @[disassembler.scala 124:19]
  wire  _T_104; // @[disassembler.scala 124:23]
  wire [7:0] Preamble01; // @[disassembler.scala 124:31]
  wire  _T_105; // @[disassembler.scala 132:16]
  wire  _T_106; // @[disassembler.scala 132:36]
  wire  _T_107; // @[disassembler.scala 132:25]
  wire [7:0] _GEN_5; // @[disassembler.scala 132:49]
  wire  _T_109; // @[disassembler.scala 152:24]
  wire  _T_110; // @[disassembler.scala 152:24]
  wire  _T_111; // @[disassembler.scala 152:24]
  wire  _T_112; // @[disassembler.scala 152:24]
  wire  _T_113; // @[disassembler.scala 152:24]
  wire  _T_114; // @[disassembler.scala 152:24]
  wire  _T_115; // @[disassembler.scala 152:24]
  wire  _T_116; // @[disassembler.scala 152:24]
  wire [2:0] _GEN_6; // @[disassembler.scala 174:37]
  wire  _T_348; // @[disassembler.scala 355:16]
  wire  _T_349; // @[disassembler.scala 355:42]
  wire  _T_350; // @[disassembler.scala 355:31]
  wire  _T_351; // @[disassembler.scala 355:69]
  wire  _T_352; // @[disassembler.scala 355:58]
  wire  DEWHITE_Result_w; // @[disassembler.scala 110:30]
  wire  _T_356; // @[disassembler.scala 358:28]
  wire  _GEN_99; // @[disassembler.scala 359:32]
  wire  _GEN_107; // @[disassembler.scala 361:32]
  wire  _GEN_115; // @[disassembler.scala 358:35]
  wire  _GEN_123; // @[disassembler.scala 356:34]
  wire  _T_375; // @[disassembler.scala 374:25]
  wire  _GEN_132; // @[disassembler.scala 374:32]
  wire  _GEN_140; // @[disassembler.scala 365:34]
  wire  _T_403; // @[disassembler.scala 381:22]
  wire  _T_407; // @[disassembler.scala 384:32]
  wire  _GEN_163; // @[disassembler.scala 384:39]
  wire  _GEN_171; // @[disassembler.scala 382:34]
  wire  _GEN_179; // @[disassembler.scala 381:29]
  wire  _GEN_188; // @[disassembler.scala 364:35]
  wire  data_w_1; // @[disassembler.scala 355:77]
  wire  _GEN_98; // @[disassembler.scala 359:32]
  wire  _GEN_106; // @[disassembler.scala 361:32]
  wire  _GEN_114; // @[disassembler.scala 358:35]
  wire  _GEN_122; // @[disassembler.scala 356:34]
  wire  _T_370; // @[disassembler.scala 374:25]
  wire  _GEN_131; // @[disassembler.scala 374:32]
  wire  _GEN_139; // @[disassembler.scala 365:34]
  wire  _GEN_162; // @[disassembler.scala 384:39]
  wire  _GEN_170; // @[disassembler.scala 382:34]
  wire  _GEN_178; // @[disassembler.scala 381:29]
  wire  _GEN_187; // @[disassembler.scala 364:35]
  wire  data_w_0; // @[disassembler.scala 355:77]
  wire [1:0] _T_127; // @[disassembler.scala 180:17]
  wire  _GEN_101; // @[disassembler.scala 359:32]
  wire  _GEN_109; // @[disassembler.scala 361:32]
  wire  _GEN_117; // @[disassembler.scala 358:35]
  wire  _GEN_125; // @[disassembler.scala 356:34]
  wire  _T_385; // @[disassembler.scala 374:25]
  wire  _GEN_134; // @[disassembler.scala 374:32]
  wire  _GEN_142; // @[disassembler.scala 365:34]
  wire  _GEN_165; // @[disassembler.scala 384:39]
  wire  _GEN_173; // @[disassembler.scala 382:34]
  wire  _GEN_181; // @[disassembler.scala 381:29]
  wire  _GEN_190; // @[disassembler.scala 364:35]
  wire  data_w_3; // @[disassembler.scala 355:77]
  wire  _GEN_100; // @[disassembler.scala 359:32]
  wire  _GEN_108; // @[disassembler.scala 361:32]
  wire  _GEN_116; // @[disassembler.scala 358:35]
  wire  _GEN_124; // @[disassembler.scala 356:34]
  wire  _T_380; // @[disassembler.scala 374:25]
  wire  _GEN_133; // @[disassembler.scala 374:32]
  wire  _GEN_141; // @[disassembler.scala 365:34]
  wire  _GEN_164; // @[disassembler.scala 384:39]
  wire  _GEN_172; // @[disassembler.scala 382:34]
  wire  _GEN_180; // @[disassembler.scala 381:29]
  wire  _GEN_189; // @[disassembler.scala 364:35]
  wire  data_w_2; // @[disassembler.scala 355:77]
  wire [1:0] _T_128; // @[disassembler.scala 180:17]
  wire [3:0] _T_129; // @[disassembler.scala 180:17]
  wire  _GEN_103; // @[disassembler.scala 359:32]
  wire  _GEN_111; // @[disassembler.scala 361:32]
  wire  _GEN_119; // @[disassembler.scala 358:35]
  wire  _GEN_127; // @[disassembler.scala 356:34]
  wire  _T_395; // @[disassembler.scala 374:25]
  wire  _GEN_136; // @[disassembler.scala 374:32]
  wire  _GEN_144; // @[disassembler.scala 365:34]
  wire  _GEN_167; // @[disassembler.scala 384:39]
  wire  _GEN_175; // @[disassembler.scala 382:34]
  wire  _GEN_183; // @[disassembler.scala 381:29]
  wire  _GEN_192; // @[disassembler.scala 364:35]
  wire  data_w_5; // @[disassembler.scala 355:77]
  wire  _GEN_102; // @[disassembler.scala 359:32]
  wire  _GEN_110; // @[disassembler.scala 361:32]
  wire  _GEN_118; // @[disassembler.scala 358:35]
  wire  _GEN_126; // @[disassembler.scala 356:34]
  wire  _T_390; // @[disassembler.scala 374:25]
  wire  _GEN_135; // @[disassembler.scala 374:32]
  wire  _GEN_143; // @[disassembler.scala 365:34]
  wire  _GEN_166; // @[disassembler.scala 384:39]
  wire  _GEN_174; // @[disassembler.scala 382:34]
  wire  _GEN_182; // @[disassembler.scala 381:29]
  wire  _GEN_191; // @[disassembler.scala 364:35]
  wire  data_w_4; // @[disassembler.scala 355:77]
  wire [1:0] _T_130; // @[disassembler.scala 180:17]
  wire  _GEN_105; // @[disassembler.scala 359:32]
  wire  _GEN_113; // @[disassembler.scala 361:32]
  wire  _GEN_121; // @[disassembler.scala 358:35]
  wire  _GEN_129; // @[disassembler.scala 356:34]
  wire  _GEN_130; // @[disassembler.scala 367:39]
  wire  _GEN_138; // @[disassembler.scala 365:34]
  wire  _GEN_169; // @[disassembler.scala 384:39]
  wire  _GEN_177; // @[disassembler.scala 382:34]
  wire  _GEN_185; // @[disassembler.scala 381:29]
  wire  _GEN_186; // @[disassembler.scala 364:35]
  wire  data_w_7; // @[disassembler.scala 355:77]
  wire  _GEN_104; // @[disassembler.scala 359:32]
  wire  _GEN_112; // @[disassembler.scala 361:32]
  wire  _GEN_120; // @[disassembler.scala 358:35]
  wire  _GEN_128; // @[disassembler.scala 356:34]
  wire  _T_400; // @[disassembler.scala 374:25]
  wire  _GEN_137; // @[disassembler.scala 374:32]
  wire  _GEN_145; // @[disassembler.scala 365:34]
  wire  _GEN_168; // @[disassembler.scala 384:39]
  wire  _GEN_176; // @[disassembler.scala 382:34]
  wire  _GEN_184; // @[disassembler.scala 381:29]
  wire  _GEN_193; // @[disassembler.scala 364:35]
  wire  data_w_6; // @[disassembler.scala 355:77]
  wire [1:0] _T_131; // @[disassembler.scala 180:17]
  wire [3:0] _T_132; // @[disassembler.scala 180:17]
  wire [7:0] _T_133; // @[disassembler.scala 180:17]
  wire  _T_134; // @[disassembler.scala 180:24]
  wire [2:0] _GEN_7; // @[disassembler.scala 180:39]
  wire [7:0] _GEN_8; // @[disassembler.scala 180:39]
  wire [2:0] _GEN_9; // @[disassembler.scala 180:39]
  wire  _T_139; // @[disassembler.scala 188:20]
  wire  _T_142; // @[disassembler.scala 188:28]
  wire [8:0] _T_148; // @[disassembler.scala 195:31]
  wire [7:0] _T_149; // @[disassembler.scala 195:31]
  wire [7:0] _GEN_10; // @[disassembler.scala 194:39]
  wire  _T_153; // @[disassembler.scala 198:29]
  wire [3:0] _T_156; // @[disassembler.scala 201:43]
  wire [2:0] _T_157; // @[disassembler.scala 201:43]
  wire [2:0] _GEN_11; // @[disassembler.scala 198:37]
  wire [2:0] _GEN_12; // @[disassembler.scala 197:36]
  wire [2:0] _GEN_13; // @[disassembler.scala 188:58]
  wire [7:0] _GEN_14; // @[disassembler.scala 188:58]
  wire [2:0] _GEN_15; // @[disassembler.scala 188:58]
  wire  _T_160; // @[disassembler.scala 206:20]
  wire  _T_163; // @[disassembler.scala 206:28]
  wire [2:0] _GEN_19; // @[disassembler.scala 206:58]
  wire [7:0] _GEN_20; // @[disassembler.scala 206:58]
  wire [2:0] _GEN_21; // @[disassembler.scala 206:58]
  wire [8:0] _T_181; // @[disassembler.scala 224:36]
  wire [8:0] _T_182; // @[disassembler.scala 224:36]
  wire [7:0] _T_183; // @[disassembler.scala 224:36]
  wire  _T_184; // @[disassembler.scala 224:20]
  wire  _T_187; // @[disassembler.scala 224:41]
  wire [2:0] _GEN_25; // @[disassembler.scala 224:71]
  wire [7:0] _GEN_26; // @[disassembler.scala 224:71]
  wire [2:0] _GEN_27; // @[disassembler.scala 224:71]
  wire  _T_205; // @[disassembler.scala 242:20]
  wire  _T_208; // @[disassembler.scala 242:28]
  wire [2:0] _GEN_31; // @[disassembler.scala 242:58]
  wire [7:0] _GEN_32; // @[disassembler.scala 242:58]
  wire [2:0] _GEN_33; // @[disassembler.scala 242:58]
  wire  _T_224; // @[disassembler.scala 259:22]
  wire  _T_229; // @[disassembler.scala 260:44]
  wire  _T_232; // @[disassembler.scala 260:81]
  wire [2:0] _GEN_34; // @[disassembler.scala 260:120]
  wire [2:0] _GEN_35; // @[disassembler.scala 259:36]
  wire [2:0] _GEN_36; // @[disassembler.scala 241:30]
  wire [7:0] _GEN_37; // @[disassembler.scala 241:30]
  wire [2:0] _GEN_38; // @[disassembler.scala 241:30]
  wire [2:0] _GEN_39; // @[disassembler.scala 223:38]
  wire [7:0] _GEN_40; // @[disassembler.scala 223:38]
  wire [2:0] _GEN_41; // @[disassembler.scala 223:38]
  wire [2:0] _GEN_42; // @[disassembler.scala 205:37]
  wire [7:0] _GEN_43; // @[disassembler.scala 205:37]
  wire [2:0] _GEN_44; // @[disassembler.scala 205:37]
  wire [2:0] _GEN_45; // @[disassembler.scala 187:29]
  wire [7:0] _GEN_46; // @[disassembler.scala 187:29]
  wire [2:0] _GEN_47; // @[disassembler.scala 187:29]
  wire [2:0] _GEN_48; // @[disassembler.scala 179:35]
  wire [7:0] _GEN_49; // @[disassembler.scala 179:35]
  wire [2:0] _GEN_50; // @[disassembler.scala 179:35]
  wire [7:0] _GEN_51; // @[disassembler.scala 167:25]
  wire  _GEN_52; // @[disassembler.scala 167:25]
  wire  _GEN_53; // @[disassembler.scala 167:25]
  wire  _GEN_54; // @[disassembler.scala 167:25]
  wire  _GEN_55; // @[disassembler.scala 167:25]
  wire  _GEN_56; // @[disassembler.scala 167:25]
  wire [2:0] state_w; // @[disassembler.scala 167:25]
  wire [7:0] counter_w; // @[disassembler.scala 167:25]
  wire [2:0] counter_byte_w; // @[disassembler.scala 167:25]
  wire  _T_236; // @[disassembler.scala 271:31]
  wire  _T_239; // @[disassembler.scala 271:52]
  wire  _T_241; // @[disassembler.scala 274:22]
  wire  _GEN_60; // @[disassembler.scala 274:32]
  wire [7:0] _GEN_61; // @[disassembler.scala 271:82]
  wire  _GEN_62; // @[disassembler.scala 271:82]
  wire  _T_245; // @[disassembler.scala 281:36]
  wire  _T_246; // @[disassembler.scala 281:23]
  wire  _T_249; // @[disassembler.scala 281:44]
  wire [7:0] _T_250; // @[disassembler.scala 282:32]
  wire  _T_251; // @[disassembler.scala 282:17]
  wire  _GEN_63; // @[disassembler.scala 282:38]
  wire  _GEN_64; // @[disassembler.scala 282:38]
  wire  _T_257; // @[disassembler.scala 286:29]
  wire  _T_260; // @[disassembler.scala 286:50]
  wire [7:0] _T_261; // @[disassembler.scala 287:32]
  wire  _T_262; // @[disassembler.scala 287:17]
  wire  _GEN_65; // @[disassembler.scala 287:39]
  wire  _GEN_66; // @[disassembler.scala 287:39]
  wire  _T_268; // @[disassembler.scala 291:29]
  wire  _T_271; // @[disassembler.scala 291:50]
  wire [7:0] _T_272; // @[disassembler.scala 292:32]
  wire  _T_273; // @[disassembler.scala 292:17]
  wire  _GEN_67; // @[disassembler.scala 292:40]
  wire  _GEN_68; // @[disassembler.scala 292:40]
  wire  _T_279; // @[disassembler.scala 296:29]
  wire  _T_282; // @[disassembler.scala 296:50]
  wire [7:0] _T_283; // @[disassembler.scala 297:32]
  wire  _T_284; // @[disassembler.scala 297:17]
  wire  _GEN_69; // @[disassembler.scala 297:40]
  wire  _GEN_71; // @[disassembler.scala 296:80]
  wire  _GEN_72; // @[disassembler.scala 296:80]
  wire  _GEN_73; // @[disassembler.scala 291:80]
  wire  _GEN_74; // @[disassembler.scala 291:80]
  wire  _GEN_75; // @[disassembler.scala 286:80]
  wire  _GEN_76; // @[disassembler.scala 286:80]
  wire  _GEN_77; // @[disassembler.scala 281:74]
  wire  _GEN_78; // @[disassembler.scala 281:74]
  wire  _T_291; // @[disassembler.scala 308:24]
  wire  _T_294; // @[disassembler.scala 308:45]
  wire [23:0] CRC_Result_w; // @[disassembler.scala 103:26]
  wire [7:0] _T_295; // @[disassembler.scala 309:33]
  wire  _T_296; // @[disassembler.scala 309:17]
  wire  _GEN_79; // @[disassembler.scala 309:39]
  wire  _GEN_80; // @[disassembler.scala 309:39]
  wire  _T_302; // @[disassembler.scala 313:30]
  wire  _T_305; // @[disassembler.scala 313:51]
  wire [7:0] _T_306; // @[disassembler.scala 314:33]
  wire  _T_307; // @[disassembler.scala 314:17]
  wire  _GEN_81; // @[disassembler.scala 314:40]
  wire  _GEN_82; // @[disassembler.scala 314:40]
  wire  _T_313; // @[disassembler.scala 318:30]
  wire  _T_316; // @[disassembler.scala 318:51]
  wire [7:0] _T_317; // @[disassembler.scala 319:33]
  wire  _T_318; // @[disassembler.scala 319:17]
  wire  _GEN_83; // @[disassembler.scala 319:41]
  wire  _GEN_85; // @[disassembler.scala 318:81]
  wire  _GEN_86; // @[disassembler.scala 318:81]
  wire  _GEN_87; // @[disassembler.scala 313:81]
  wire  _GEN_88; // @[disassembler.scala 313:81]
  wire  _GEN_89; // @[disassembler.scala 308:75]
  wire  _GEN_90; // @[disassembler.scala 308:75]
  wire  _T_330; // @[disassembler.scala 334:33]
  wire  _GEN_91; // @[disassembler.scala 336:43]
  wire  _GEN_92; // @[disassembler.scala 334:60]
  wire  _GEN_93; // @[disassembler.scala 331:49]
  wire  _GEN_94; // @[disassembler.scala 349:43]
  wire  _GEN_95; // @[disassembler.scala 347:60]
  wire  _GEN_96; // @[disassembler.scala 344:35]
  wire  _GEN_97; // @[disassembler.scala 342:25]
  wire  CRC_Data_w; // @[disassembler.scala 396:58]
  wire  CRC_Valid_w; // @[disassembler.scala 396:58]
  wire  DEWHITE_Data_w; // @[disassembler.scala 408:77]
  wire  DEWHITE_Valid_w; // @[disassembler.scala 408:77]
  ble_crc CRC_inst ( // @[disassembler.scala 425:24]
    .clock(CRC_inst_clock),
    .reset(CRC_inst_reset),
    .io_operand_valid(CRC_inst_io_operand_valid),
    .io_operand_bits(CRC_inst_io_operand_bits),
    .io_result_bits(CRC_inst_io_result_bits),
    .io_seed(CRC_inst_io_seed),
    .io_init(CRC_inst_io_init)
  );
  ble_whitening WHITE_inst ( // @[disassembler.scala 435:26]
    .clock(WHITE_inst_clock),
    .reset(WHITE_inst_reset),
    .io_operand_valid(WHITE_inst_io_operand_valid),
    .io_operand_bits(WHITE_inst_io_operand_bits),
    .io_result_bits(WHITE_inst_io_result_bits),
    .io_seed(WHITE_inst_io_seed),
    .io_init(WHITE_inst_io_init)
  );
  assign DMA_Data_Fire_w = io_DMA_Data_o_ready & io_DMA_Data_o_valid; // @[disassembler.scala 115:42]
  assign AFIFO_Fire_w = io_AFIFO_Data_i_ready & io_AFIFO_Data_i_valid; // @[disassembler.scala 116:41]
  assign _T_102 = io_REG_AA_i[0]; // @[disassembler.scala 124:19]
  assign _T_104 = _T_102 == 1'h0; // @[disassembler.scala 124:23]
  assign Preamble01 = _T_104 ? 8'haa : 8'h55; // @[disassembler.scala 124:31]
  assign _T_105 = state_r == 3'h0; // @[disassembler.scala 132:16]
  assign _T_106 = state_r == 3'h1; // @[disassembler.scala 132:36]
  assign _T_107 = _T_105 | _T_106; // @[disassembler.scala 132:25]
  assign _GEN_5 = _T_107 ? 8'h0 : data_r; // @[disassembler.scala 132:49]
  assign _T_109 = data_r[0]; // @[disassembler.scala 152:24]
  assign _T_110 = data_r[1]; // @[disassembler.scala 152:24]
  assign _T_111 = data_r[2]; // @[disassembler.scala 152:24]
  assign _T_112 = data_r[3]; // @[disassembler.scala 152:24]
  assign _T_113 = data_r[4]; // @[disassembler.scala 152:24]
  assign _T_114 = data_r[5]; // @[disassembler.scala 152:24]
  assign _T_115 = data_r[6]; // @[disassembler.scala 152:24]
  assign _T_116 = data_r[7]; // @[disassembler.scala 152:24]
  assign _GEN_6 = io_DMA_Switch_i ? 3'h1 : 3'h0; // @[disassembler.scala 174:37]
  assign _T_348 = state_r == 3'h3; // @[disassembler.scala 355:16]
  assign _T_349 = state_r == 3'h4; // @[disassembler.scala 355:42]
  assign _T_350 = _T_348 | _T_349; // @[disassembler.scala 355:31]
  assign _T_351 = state_r == 3'h5; // @[disassembler.scala 355:69]
  assign _T_352 = _T_350 | _T_351; // @[disassembler.scala 355:58]
  assign DEWHITE_Result_w = WHITE_inst_io_result_bits; // @[disassembler.scala 110:30]
  assign _T_356 = DEWHITE_Result_w == 1'h0; // @[disassembler.scala 358:28]
  assign _GEN_99 = 3'h1 == counter_byte_r ? 1'h0 : _T_110; // @[disassembler.scala 359:32]
  assign _GEN_107 = 3'h1 == counter_byte_r ? 1'h1 : _T_110; // @[disassembler.scala 361:32]
  assign _GEN_115 = _T_356 ? _GEN_99 : _GEN_107; // @[disassembler.scala 358:35]
  assign _GEN_123 = AFIFO_Fire_w ? _GEN_115 : _T_110; // @[disassembler.scala 356:34]
  assign _T_375 = _T_111 == 1'h0; // @[disassembler.scala 374:25]
  assign _GEN_132 = _T_375 ? 1'h0 : 1'h1; // @[disassembler.scala 374:32]
  assign _GEN_140 = AFIFO_Fire_w ? _GEN_132 : _T_110; // @[disassembler.scala 365:34]
  assign _T_403 = state_r == 3'h2; // @[disassembler.scala 381:22]
  assign _T_407 = io_AFIFO_Data_i_bits == 1'h0; // @[disassembler.scala 384:32]
  assign _GEN_163 = _T_407 ? _GEN_99 : _GEN_107; // @[disassembler.scala 384:39]
  assign _GEN_171 = AFIFO_Fire_w ? _GEN_163 : _T_110; // @[disassembler.scala 382:34]
  assign _GEN_179 = _T_403 ? _GEN_171 : _T_110; // @[disassembler.scala 381:29]
  assign _GEN_188 = _T_106 ? _GEN_140 : _GEN_179; // @[disassembler.scala 364:35]
  assign data_w_1 = _T_352 ? _GEN_123 : _GEN_188; // @[disassembler.scala 355:77]
  assign _GEN_98 = 3'h0 == counter_byte_r ? 1'h0 : _T_109; // @[disassembler.scala 359:32]
  assign _GEN_106 = 3'h0 == counter_byte_r ? 1'h1 : _T_109; // @[disassembler.scala 361:32]
  assign _GEN_114 = _T_356 ? _GEN_98 : _GEN_106; // @[disassembler.scala 358:35]
  assign _GEN_122 = AFIFO_Fire_w ? _GEN_114 : _T_109; // @[disassembler.scala 356:34]
  assign _T_370 = _T_110 == 1'h0; // @[disassembler.scala 374:25]
  assign _GEN_131 = _T_370 ? 1'h0 : 1'h1; // @[disassembler.scala 374:32]
  assign _GEN_139 = AFIFO_Fire_w ? _GEN_131 : _T_109; // @[disassembler.scala 365:34]
  assign _GEN_162 = _T_407 ? _GEN_98 : _GEN_106; // @[disassembler.scala 384:39]
  assign _GEN_170 = AFIFO_Fire_w ? _GEN_162 : _T_109; // @[disassembler.scala 382:34]
  assign _GEN_178 = _T_403 ? _GEN_170 : _T_109; // @[disassembler.scala 381:29]
  assign _GEN_187 = _T_106 ? _GEN_139 : _GEN_178; // @[disassembler.scala 364:35]
  assign data_w_0 = _T_352 ? _GEN_122 : _GEN_187; // @[disassembler.scala 355:77]
  assign _T_127 = {data_w_1,data_w_0}; // @[disassembler.scala 180:17]
  assign _GEN_101 = 3'h3 == counter_byte_r ? 1'h0 : _T_112; // @[disassembler.scala 359:32]
  assign _GEN_109 = 3'h3 == counter_byte_r ? 1'h1 : _T_112; // @[disassembler.scala 361:32]
  assign _GEN_117 = _T_356 ? _GEN_101 : _GEN_109; // @[disassembler.scala 358:35]
  assign _GEN_125 = AFIFO_Fire_w ? _GEN_117 : _T_112; // @[disassembler.scala 356:34]
  assign _T_385 = _T_113 == 1'h0; // @[disassembler.scala 374:25]
  assign _GEN_134 = _T_385 ? 1'h0 : 1'h1; // @[disassembler.scala 374:32]
  assign _GEN_142 = AFIFO_Fire_w ? _GEN_134 : _T_112; // @[disassembler.scala 365:34]
  assign _GEN_165 = _T_407 ? _GEN_101 : _GEN_109; // @[disassembler.scala 384:39]
  assign _GEN_173 = AFIFO_Fire_w ? _GEN_165 : _T_112; // @[disassembler.scala 382:34]
  assign _GEN_181 = _T_403 ? _GEN_173 : _T_112; // @[disassembler.scala 381:29]
  assign _GEN_190 = _T_106 ? _GEN_142 : _GEN_181; // @[disassembler.scala 364:35]
  assign data_w_3 = _T_352 ? _GEN_125 : _GEN_190; // @[disassembler.scala 355:77]
  assign _GEN_100 = 3'h2 == counter_byte_r ? 1'h0 : _T_111; // @[disassembler.scala 359:32]
  assign _GEN_108 = 3'h2 == counter_byte_r ? 1'h1 : _T_111; // @[disassembler.scala 361:32]
  assign _GEN_116 = _T_356 ? _GEN_100 : _GEN_108; // @[disassembler.scala 358:35]
  assign _GEN_124 = AFIFO_Fire_w ? _GEN_116 : _T_111; // @[disassembler.scala 356:34]
  assign _T_380 = _T_112 == 1'h0; // @[disassembler.scala 374:25]
  assign _GEN_133 = _T_380 ? 1'h0 : 1'h1; // @[disassembler.scala 374:32]
  assign _GEN_141 = AFIFO_Fire_w ? _GEN_133 : _T_111; // @[disassembler.scala 365:34]
  assign _GEN_164 = _T_407 ? _GEN_100 : _GEN_108; // @[disassembler.scala 384:39]
  assign _GEN_172 = AFIFO_Fire_w ? _GEN_164 : _T_111; // @[disassembler.scala 382:34]
  assign _GEN_180 = _T_403 ? _GEN_172 : _T_111; // @[disassembler.scala 381:29]
  assign _GEN_189 = _T_106 ? _GEN_141 : _GEN_180; // @[disassembler.scala 364:35]
  assign data_w_2 = _T_352 ? _GEN_124 : _GEN_189; // @[disassembler.scala 355:77]
  assign _T_128 = {data_w_3,data_w_2}; // @[disassembler.scala 180:17]
  assign _T_129 = {_T_128,_T_127}; // @[disassembler.scala 180:17]
  assign _GEN_103 = 3'h5 == counter_byte_r ? 1'h0 : _T_114; // @[disassembler.scala 359:32]
  assign _GEN_111 = 3'h5 == counter_byte_r ? 1'h1 : _T_114; // @[disassembler.scala 361:32]
  assign _GEN_119 = _T_356 ? _GEN_103 : _GEN_111; // @[disassembler.scala 358:35]
  assign _GEN_127 = AFIFO_Fire_w ? _GEN_119 : _T_114; // @[disassembler.scala 356:34]
  assign _T_395 = _T_115 == 1'h0; // @[disassembler.scala 374:25]
  assign _GEN_136 = _T_395 ? 1'h0 : 1'h1; // @[disassembler.scala 374:32]
  assign _GEN_144 = AFIFO_Fire_w ? _GEN_136 : _T_114; // @[disassembler.scala 365:34]
  assign _GEN_167 = _T_407 ? _GEN_103 : _GEN_111; // @[disassembler.scala 384:39]
  assign _GEN_175 = AFIFO_Fire_w ? _GEN_167 : _T_114; // @[disassembler.scala 382:34]
  assign _GEN_183 = _T_403 ? _GEN_175 : _T_114; // @[disassembler.scala 381:29]
  assign _GEN_192 = _T_106 ? _GEN_144 : _GEN_183; // @[disassembler.scala 364:35]
  assign data_w_5 = _T_352 ? _GEN_127 : _GEN_192; // @[disassembler.scala 355:77]
  assign _GEN_102 = 3'h4 == counter_byte_r ? 1'h0 : _T_113; // @[disassembler.scala 359:32]
  assign _GEN_110 = 3'h4 == counter_byte_r ? 1'h1 : _T_113; // @[disassembler.scala 361:32]
  assign _GEN_118 = _T_356 ? _GEN_102 : _GEN_110; // @[disassembler.scala 358:35]
  assign _GEN_126 = AFIFO_Fire_w ? _GEN_118 : _T_113; // @[disassembler.scala 356:34]
  assign _T_390 = _T_114 == 1'h0; // @[disassembler.scala 374:25]
  assign _GEN_135 = _T_390 ? 1'h0 : 1'h1; // @[disassembler.scala 374:32]
  assign _GEN_143 = AFIFO_Fire_w ? _GEN_135 : _T_113; // @[disassembler.scala 365:34]
  assign _GEN_166 = _T_407 ? _GEN_102 : _GEN_110; // @[disassembler.scala 384:39]
  assign _GEN_174 = AFIFO_Fire_w ? _GEN_166 : _T_113; // @[disassembler.scala 382:34]
  assign _GEN_182 = _T_403 ? _GEN_174 : _T_113; // @[disassembler.scala 381:29]
  assign _GEN_191 = _T_106 ? _GEN_143 : _GEN_182; // @[disassembler.scala 364:35]
  assign data_w_4 = _T_352 ? _GEN_126 : _GEN_191; // @[disassembler.scala 355:77]
  assign _T_130 = {data_w_5,data_w_4}; // @[disassembler.scala 180:17]
  assign _GEN_105 = 3'h7 == counter_byte_r ? 1'h0 : _T_116; // @[disassembler.scala 359:32]
  assign _GEN_113 = 3'h7 == counter_byte_r ? 1'h1 : _T_116; // @[disassembler.scala 361:32]
  assign _GEN_121 = _T_356 ? _GEN_105 : _GEN_113; // @[disassembler.scala 358:35]
  assign _GEN_129 = AFIFO_Fire_w ? _GEN_121 : _T_116; // @[disassembler.scala 356:34]
  assign _GEN_130 = _T_407 ? 1'h0 : 1'h1; // @[disassembler.scala 367:39]
  assign _GEN_138 = AFIFO_Fire_w ? _GEN_130 : _T_116; // @[disassembler.scala 365:34]
  assign _GEN_169 = _T_407 ? _GEN_105 : _GEN_113; // @[disassembler.scala 384:39]
  assign _GEN_177 = AFIFO_Fire_w ? _GEN_169 : _T_116; // @[disassembler.scala 382:34]
  assign _GEN_185 = _T_403 ? _GEN_177 : _T_116; // @[disassembler.scala 381:29]
  assign _GEN_186 = _T_106 ? _GEN_138 : _GEN_185; // @[disassembler.scala 364:35]
  assign data_w_7 = _T_352 ? _GEN_129 : _GEN_186; // @[disassembler.scala 355:77]
  assign _GEN_104 = 3'h6 == counter_byte_r ? 1'h0 : _T_115; // @[disassembler.scala 359:32]
  assign _GEN_112 = 3'h6 == counter_byte_r ? 1'h1 : _T_115; // @[disassembler.scala 361:32]
  assign _GEN_120 = _T_356 ? _GEN_104 : _GEN_112; // @[disassembler.scala 358:35]
  assign _GEN_128 = AFIFO_Fire_w ? _GEN_120 : _T_115; // @[disassembler.scala 356:34]
  assign _T_400 = _T_116 == 1'h0; // @[disassembler.scala 374:25]
  assign _GEN_137 = _T_400 ? 1'h0 : 1'h1; // @[disassembler.scala 374:32]
  assign _GEN_145 = AFIFO_Fire_w ? _GEN_137 : _T_115; // @[disassembler.scala 365:34]
  assign _GEN_168 = _T_407 ? _GEN_104 : _GEN_112; // @[disassembler.scala 384:39]
  assign _GEN_176 = AFIFO_Fire_w ? _GEN_168 : _T_115; // @[disassembler.scala 382:34]
  assign _GEN_184 = _T_403 ? _GEN_176 : _T_115; // @[disassembler.scala 381:29]
  assign _GEN_193 = _T_106 ? _GEN_145 : _GEN_184; // @[disassembler.scala 364:35]
  assign data_w_6 = _T_352 ? _GEN_128 : _GEN_193; // @[disassembler.scala 355:77]
  assign _T_131 = {data_w_7,data_w_6}; // @[disassembler.scala 180:17]
  assign _T_132 = {_T_131,_T_130}; // @[disassembler.scala 180:17]
  assign _T_133 = {_T_132,_T_129}; // @[disassembler.scala 180:17]
  assign _T_134 = _T_133 == Preamble01; // @[disassembler.scala 180:24]
  assign _GEN_7 = _T_134 ? 3'h2 : 3'h1; // @[disassembler.scala 180:39]
  assign _GEN_8 = _T_134 ? 8'h0 : counter_r; // @[disassembler.scala 180:39]
  assign _GEN_9 = _T_134 ? 3'h0 : counter_byte_r; // @[disassembler.scala 180:39]
  assign _T_139 = counter_r == 8'h3; // @[disassembler.scala 188:20]
  assign _T_142 = _T_139 & DMA_Data_Fire_w; // @[disassembler.scala 188:28]
  assign _T_148 = counter_r + 8'h1; // @[disassembler.scala 195:31]
  assign _T_149 = _T_148[7:0]; // @[disassembler.scala 195:31]
  assign _GEN_10 = DMA_Data_Fire_w ? _T_149 : counter_r; // @[disassembler.scala 194:39]
  assign _T_153 = counter_byte_r == 3'h7; // @[disassembler.scala 198:29]
  assign _T_156 = counter_byte_r + 3'h1; // @[disassembler.scala 201:43]
  assign _T_157 = _T_156[2:0]; // @[disassembler.scala 201:43]
  assign _GEN_11 = _T_153 ? 3'h0 : _T_157; // @[disassembler.scala 198:37]
  assign _GEN_12 = AFIFO_Fire_w ? _GEN_11 : counter_byte_r; // @[disassembler.scala 197:36]
  assign _GEN_13 = _T_142 ? 3'h3 : 3'h2; // @[disassembler.scala 188:58]
  assign _GEN_14 = _T_142 ? 8'h0 : _GEN_10; // @[disassembler.scala 188:58]
  assign _GEN_15 = _T_142 ? 3'h0 : _GEN_12; // @[disassembler.scala 188:58]
  assign _T_160 = counter_r == 8'h1; // @[disassembler.scala 206:20]
  assign _T_163 = _T_160 & DMA_Data_Fire_w; // @[disassembler.scala 206:28]
  assign _GEN_19 = _T_163 ? 3'h4 : 3'h3; // @[disassembler.scala 206:58]
  assign _GEN_20 = _T_163 ? 8'h0 : _GEN_10; // @[disassembler.scala 206:58]
  assign _GEN_21 = _T_163 ? 3'h0 : _GEN_12; // @[disassembler.scala 206:58]
  assign _T_181 = PDU_Length_r - 8'h1; // @[disassembler.scala 224:36]
  assign _T_182 = $unsigned(_T_181); // @[disassembler.scala 224:36]
  assign _T_183 = _T_182[7:0]; // @[disassembler.scala 224:36]
  assign _T_184 = counter_r == _T_183; // @[disassembler.scala 224:20]
  assign _T_187 = _T_184 & DMA_Data_Fire_w; // @[disassembler.scala 224:41]
  assign _GEN_25 = _T_187 ? 3'h5 : 3'h4; // @[disassembler.scala 224:71]
  assign _GEN_26 = _T_187 ? 8'h0 : _GEN_10; // @[disassembler.scala 224:71]
  assign _GEN_27 = _T_187 ? 3'h0 : _GEN_12; // @[disassembler.scala 224:71]
  assign _T_205 = counter_r == 8'h2; // @[disassembler.scala 242:20]
  assign _T_208 = _T_205 & DMA_Data_Fire_w; // @[disassembler.scala 242:28]
  assign _GEN_31 = _T_208 ? 3'h6 : 3'h5; // @[disassembler.scala 242:58]
  assign _GEN_32 = _T_208 ? 8'h0 : _GEN_10; // @[disassembler.scala 242:58]
  assign _GEN_33 = _T_208 ? 3'h0 : _GEN_12; // @[disassembler.scala 242:58]
  assign _T_224 = state_r == 3'h6; // @[disassembler.scala 259:22]
  assign _T_229 = io_DMA_Length_o_ready & io_DMA_Flag_AA_o_ready; // @[disassembler.scala 260:44]
  assign _T_232 = _T_229 & io_DMA_Flag_CRC_o_ready; // @[disassembler.scala 260:81]
  assign _GEN_34 = _T_232 ? 3'h0 : 3'h6; // @[disassembler.scala 260:120]
  assign _GEN_35 = _T_224 ? _GEN_34 : 3'h0; // @[disassembler.scala 259:36]
  assign _GEN_36 = _T_351 ? _GEN_31 : _GEN_35; // @[disassembler.scala 241:30]
  assign _GEN_37 = _T_351 ? _GEN_32 : counter_r; // @[disassembler.scala 241:30]
  assign _GEN_38 = _T_351 ? _GEN_33 : counter_byte_r; // @[disassembler.scala 241:30]
  assign _GEN_39 = _T_349 ? _GEN_25 : _GEN_36; // @[disassembler.scala 223:38]
  assign _GEN_40 = _T_349 ? _GEN_26 : _GEN_37; // @[disassembler.scala 223:38]
  assign _GEN_41 = _T_349 ? _GEN_27 : _GEN_38; // @[disassembler.scala 223:38]
  assign _GEN_42 = _T_348 ? _GEN_19 : _GEN_39; // @[disassembler.scala 205:37]
  assign _GEN_43 = _T_348 ? _GEN_20 : _GEN_40; // @[disassembler.scala 205:37]
  assign _GEN_44 = _T_348 ? _GEN_21 : _GEN_41; // @[disassembler.scala 205:37]
  assign _GEN_45 = _T_403 ? _GEN_13 : _GEN_42; // @[disassembler.scala 187:29]
  assign _GEN_46 = _T_403 ? _GEN_14 : _GEN_43; // @[disassembler.scala 187:29]
  assign _GEN_47 = _T_403 ? _GEN_15 : _GEN_44; // @[disassembler.scala 187:29]
  assign _GEN_48 = _T_106 ? _GEN_7 : _GEN_45; // @[disassembler.scala 179:35]
  assign _GEN_49 = _T_106 ? _GEN_8 : _GEN_46; // @[disassembler.scala 179:35]
  assign _GEN_50 = _T_106 ? _GEN_9 : _GEN_47; // @[disassembler.scala 179:35]
  assign _GEN_51 = _T_105 ? 8'h0 : PDU_Length_r; // @[disassembler.scala 167:25]
  assign _GEN_52 = _T_105 ? 1'h0 : PDU_Length_Valid_r; // @[disassembler.scala 167:25]
  assign _GEN_53 = _T_105 ? 1'h0 : Flag_AA_r; // @[disassembler.scala 167:25]
  assign _GEN_54 = _T_105 ? 1'h0 : Flag_AA_Valid_r; // @[disassembler.scala 167:25]
  assign _GEN_55 = _T_105 ? 1'h0 : Flag_CRC_r; // @[disassembler.scala 167:25]
  assign _GEN_56 = _T_105 ? 1'h0 : Flag_CRC_Valid_r; // @[disassembler.scala 167:25]
  assign state_w = _T_105 ? _GEN_6 : _GEN_48; // @[disassembler.scala 167:25]
  assign counter_w = _T_105 ? counter_r : _GEN_49; // @[disassembler.scala 167:25]
  assign counter_byte_w = _T_105 ? counter_byte_r : _GEN_50; // @[disassembler.scala 167:25]
  assign _T_236 = _T_348 & _T_160; // @[disassembler.scala 271:31]
  assign _T_239 = _T_236 & DMA_Data_Fire_w; // @[disassembler.scala 271:52]
  assign _T_241 = state_w == 3'h0; // @[disassembler.scala 274:22]
  assign _GEN_60 = _T_241 ? 1'h0 : _GEN_52; // @[disassembler.scala 274:32]
  assign _GEN_61 = _T_239 ? data_r : _GEN_51; // @[disassembler.scala 271:82]
  assign _GEN_62 = _T_239 ? 1'h1 : _GEN_60; // @[disassembler.scala 271:82]
  assign _T_245 = counter_r == 8'h0; // @[disassembler.scala 281:36]
  assign _T_246 = _T_403 & _T_245; // @[disassembler.scala 281:23]
  assign _T_249 = _T_246 & DMA_Data_Fire_w; // @[disassembler.scala 281:44]
  assign _T_250 = io_REG_AA_i[7:0]; // @[disassembler.scala 282:32]
  assign _T_251 = data_r != _T_250; // @[disassembler.scala 282:17]
  assign _GEN_63 = _T_251 ? 1'h1 : _GEN_53; // @[disassembler.scala 282:38]
  assign _GEN_64 = _T_251 ? 1'h1 : _GEN_54; // @[disassembler.scala 282:38]
  assign _T_257 = _T_403 & _T_160; // @[disassembler.scala 286:29]
  assign _T_260 = _T_257 & DMA_Data_Fire_w; // @[disassembler.scala 286:50]
  assign _T_261 = io_REG_AA_i[15:8]; // @[disassembler.scala 287:32]
  assign _T_262 = data_r != _T_261; // @[disassembler.scala 287:17]
  assign _GEN_65 = _T_262 ? 1'h1 : _GEN_53; // @[disassembler.scala 287:39]
  assign _GEN_66 = _T_262 ? 1'h1 : _GEN_54; // @[disassembler.scala 287:39]
  assign _T_268 = _T_403 & _T_205; // @[disassembler.scala 291:29]
  assign _T_271 = _T_268 & DMA_Data_Fire_w; // @[disassembler.scala 291:50]
  assign _T_272 = io_REG_AA_i[23:16]; // @[disassembler.scala 292:32]
  assign _T_273 = data_r != _T_272; // @[disassembler.scala 292:17]
  assign _GEN_67 = _T_273 ? 1'h1 : _GEN_53; // @[disassembler.scala 292:40]
  assign _GEN_68 = _T_273 ? 1'h1 : _GEN_54; // @[disassembler.scala 292:40]
  assign _T_279 = _T_403 & _T_139; // @[disassembler.scala 296:29]
  assign _T_282 = _T_279 & DMA_Data_Fire_w; // @[disassembler.scala 296:50]
  assign _T_283 = io_REG_AA_i[31:24]; // @[disassembler.scala 297:32]
  assign _T_284 = data_r != _T_283; // @[disassembler.scala 297:17]
  assign _GEN_69 = _T_284 ? 1'h1 : _GEN_53; // @[disassembler.scala 297:40]
  assign _GEN_71 = _T_282 ? _GEN_69 : _GEN_53; // @[disassembler.scala 296:80]
  assign _GEN_72 = _T_282 ? 1'h1 : _GEN_54; // @[disassembler.scala 296:80]
  assign _GEN_73 = _T_271 ? _GEN_67 : _GEN_71; // @[disassembler.scala 291:80]
  assign _GEN_74 = _T_271 ? _GEN_68 : _GEN_72; // @[disassembler.scala 291:80]
  assign _GEN_75 = _T_260 ? _GEN_65 : _GEN_73; // @[disassembler.scala 286:80]
  assign _GEN_76 = _T_260 ? _GEN_66 : _GEN_74; // @[disassembler.scala 286:80]
  assign _GEN_77 = _T_249 ? _GEN_63 : _GEN_75; // @[disassembler.scala 281:74]
  assign _GEN_78 = _T_249 ? _GEN_64 : _GEN_76; // @[disassembler.scala 281:74]
  assign _T_291 = _T_351 & _T_245; // @[disassembler.scala 308:24]
  assign _T_294 = _T_291 & DMA_Data_Fire_w; // @[disassembler.scala 308:45]
  assign CRC_Result_w = CRC_inst_io_result_bits; // @[disassembler.scala 103:26]
  assign _T_295 = CRC_Result_w[7:0]; // @[disassembler.scala 309:33]
  assign _T_296 = data_r != _T_295; // @[disassembler.scala 309:17]
  assign _GEN_79 = _T_296 ? 1'h1 : _GEN_55; // @[disassembler.scala 309:39]
  assign _GEN_80 = _T_296 ? 1'h1 : _GEN_56; // @[disassembler.scala 309:39]
  assign _T_302 = _T_351 & _T_160; // @[disassembler.scala 313:30]
  assign _T_305 = _T_302 & DMA_Data_Fire_w; // @[disassembler.scala 313:51]
  assign _T_306 = CRC_Result_w[15:8]; // @[disassembler.scala 314:33]
  assign _T_307 = data_r != _T_306; // @[disassembler.scala 314:17]
  assign _GEN_81 = _T_307 ? 1'h1 : _GEN_55; // @[disassembler.scala 314:40]
  assign _GEN_82 = _T_307 ? 1'h1 : _GEN_56; // @[disassembler.scala 314:40]
  assign _T_313 = _T_351 & _T_205; // @[disassembler.scala 318:30]
  assign _T_316 = _T_313 & DMA_Data_Fire_w; // @[disassembler.scala 318:51]
  assign _T_317 = CRC_Result_w[23:16]; // @[disassembler.scala 319:33]
  assign _T_318 = data_r != _T_317; // @[disassembler.scala 319:17]
  assign _GEN_83 = _T_318 ? 1'h1 : _GEN_55; // @[disassembler.scala 319:41]
  assign _GEN_85 = _T_316 ? _GEN_83 : _GEN_55; // @[disassembler.scala 318:81]
  assign _GEN_86 = _T_316 ? 1'h1 : _GEN_56; // @[disassembler.scala 318:81]
  assign _GEN_87 = _T_305 ? _GEN_81 : _GEN_85; // @[disassembler.scala 313:81]
  assign _GEN_88 = _T_305 ? _GEN_82 : _GEN_86; // @[disassembler.scala 313:81]
  assign _GEN_89 = _T_294 ? _GEN_79 : _GEN_87; // @[disassembler.scala 308:75]
  assign _GEN_90 = _T_294 ? _GEN_80 : _GEN_88; // @[disassembler.scala 308:75]
  assign _T_330 = _T_153 & AFIFO_Fire_w; // @[disassembler.scala 334:33]
  assign _GEN_91 = DMA_Data_Fire_w ? 1'h0 : DMA_Data_Valid_r; // @[disassembler.scala 336:43]
  assign _GEN_92 = _T_330 ? 1'h1 : _GEN_91; // @[disassembler.scala 334:60]
  assign _GEN_93 = _T_107 ? 1'h0 : _GEN_92; // @[disassembler.scala 331:49]
  assign _GEN_94 = DMA_Data_Fire_w ? 1'h1 : AFIFO_Ready_r; // @[disassembler.scala 349:43]
  assign _GEN_95 = _T_330 ? 1'h0 : _GEN_94; // @[disassembler.scala 347:60]
  assign _GEN_96 = _T_106 ? 1'h1 : _GEN_95; // @[disassembler.scala 344:35]
  assign _GEN_97 = _T_105 ? 1'h0 : _GEN_96; // @[disassembler.scala 342:25]
  assign CRC_Data_w = _T_350 ? DEWHITE_Result_w : 1'h0; // @[disassembler.scala 396:58]
  assign CRC_Valid_w = _T_350 ? AFIFO_Fire_w : 1'h0; // @[disassembler.scala 396:58]
  assign DEWHITE_Data_w = _T_352 ? io_AFIFO_Data_i_bits : 1'h0; // @[disassembler.scala 408:77]
  assign DEWHITE_Valid_w = _T_352 ? AFIFO_Fire_w : 1'h0; // @[disassembler.scala 408:77]
  assign io_DMA_Data_o_valid = DMA_Data_Valid_r;
  assign io_DMA_Data_o_bits = _GEN_5;
  assign io_DMA_Length_o_valid = PDU_Length_Valid_r;
  assign io_DMA_Length_o_bits = PDU_Length_r;
  assign io_DMA_Flag_AA_o_valid = Flag_AA_Valid_r;
  assign io_DMA_Flag_AA_o_bits = Flag_AA_r;
  assign io_DMA_Flag_CRC_o_valid = Flag_CRC_Valid_r;
  assign io_DMA_Flag_CRC_o_bits = Flag_CRC_r;
  assign io_AFIFO_Data_i_ready = AFIFO_Ready_r;
  assign CRC_inst_clock = clock;
  assign CRC_inst_reset = reset;
  assign CRC_inst_io_operand_valid = CRC_Valid_w;
  assign CRC_inst_io_operand_bits = CRC_Data_w;
  assign CRC_inst_io_seed = io_REG_CRC_Seed_i;
  assign CRC_inst_io_init = _T_105;
  assign WHITE_inst_clock = clock;
  assign WHITE_inst_reset = reset;
  assign WHITE_inst_io_operand_valid = DEWHITE_Valid_w;
  assign WHITE_inst_io_operand_bits = DEWHITE_Data_w;
  assign WHITE_inst_io_seed = io_REG_DeWhite_Seed_i;
  assign WHITE_inst_io_init = _T_105;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  state_r = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  counter_r = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  counter_byte_r = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  PDU_Length_r = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  PDU_Length_Valid_r = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  Flag_AA_r = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  Flag_AA_Valid_r = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  Flag_CRC_r = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  Flag_CRC_Valid_r = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  DMA_Data_Valid_r = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  AFIFO_Ready_r = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  data_r = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state_r <= 3'h0;
    end else begin
      if (_T_105) begin
        if (io_DMA_Switch_i) begin
          state_r <= 3'h1;
        end else begin
          state_r <= 3'h0;
        end
      end else begin
        if (_T_106) begin
          if (_T_134) begin
            state_r <= 3'h2;
          end else begin
            state_r <= 3'h1;
          end
        end else begin
          if (_T_403) begin
            if (_T_142) begin
              state_r <= 3'h3;
            end else begin
              state_r <= 3'h2;
            end
          end else begin
            if (_T_348) begin
              if (_T_163) begin
                state_r <= 3'h4;
              end else begin
                state_r <= 3'h3;
              end
            end else begin
              if (_T_349) begin
                if (_T_187) begin
                  state_r <= 3'h5;
                end else begin
                  state_r <= 3'h4;
                end
              end else begin
                if (_T_351) begin
                  if (_T_208) begin
                    state_r <= 3'h6;
                  end else begin
                    state_r <= 3'h5;
                  end
                end else begin
                  if (_T_224) begin
                    if (_T_232) begin
                      state_r <= 3'h0;
                    end else begin
                      state_r <= 3'h6;
                    end
                  end else begin
                    state_r <= 3'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      counter_r <= 8'h0;
    end else begin
      if (!(_T_105)) begin
        if (_T_106) begin
          if (_T_134) begin
            counter_r <= 8'h0;
          end
        end else begin
          if (_T_403) begin
            if (_T_142) begin
              counter_r <= 8'h0;
            end else begin
              if (DMA_Data_Fire_w) begin
                counter_r <= _T_149;
              end
            end
          end else begin
            if (_T_348) begin
              if (_T_163) begin
                counter_r <= 8'h0;
              end else begin
                if (DMA_Data_Fire_w) begin
                  counter_r <= _T_149;
                end
              end
            end else begin
              if (_T_349) begin
                if (_T_187) begin
                  counter_r <= 8'h0;
                end else begin
                  if (DMA_Data_Fire_w) begin
                    counter_r <= _T_149;
                  end
                end
              end else begin
                if (_T_351) begin
                  if (_T_208) begin
                    counter_r <= 8'h0;
                  end else begin
                    if (DMA_Data_Fire_w) begin
                      counter_r <= _T_149;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      counter_byte_r <= 3'h0;
    end else begin
      if (!(_T_105)) begin
        if (_T_106) begin
          if (_T_134) begin
            counter_byte_r <= 3'h0;
          end
        end else begin
          if (_T_403) begin
            if (_T_142) begin
              counter_byte_r <= 3'h0;
            end else begin
              if (AFIFO_Fire_w) begin
                if (_T_153) begin
                  counter_byte_r <= 3'h0;
                end else begin
                  counter_byte_r <= _T_157;
                end
              end
            end
          end else begin
            if (_T_348) begin
              if (_T_163) begin
                counter_byte_r <= 3'h0;
              end else begin
                if (AFIFO_Fire_w) begin
                  if (_T_153) begin
                    counter_byte_r <= 3'h0;
                  end else begin
                    counter_byte_r <= _T_157;
                  end
                end
              end
            end else begin
              if (_T_349) begin
                if (_T_187) begin
                  counter_byte_r <= 3'h0;
                end else begin
                  if (AFIFO_Fire_w) begin
                    if (_T_153) begin
                      counter_byte_r <= 3'h0;
                    end else begin
                      counter_byte_r <= _T_157;
                    end
                  end
                end
              end else begin
                if (_T_351) begin
                  if (_T_208) begin
                    counter_byte_r <= 3'h0;
                  end else begin
                    if (AFIFO_Fire_w) begin
                      if (_T_153) begin
                        counter_byte_r <= 3'h0;
                      end else begin
                        counter_byte_r <= _T_157;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      PDU_Length_r <= 8'h0;
    end else begin
      if (_T_239) begin
        PDU_Length_r <= data_r;
      end else begin
        if (_T_105) begin
          PDU_Length_r <= 8'h0;
        end
      end
    end
    if (reset) begin
      PDU_Length_Valid_r <= 1'h0;
    end else begin
      if (_T_239) begin
        PDU_Length_Valid_r <= 1'h1;
      end else begin
        if (_T_241) begin
          PDU_Length_Valid_r <= 1'h0;
        end else begin
          if (_T_105) begin
            PDU_Length_Valid_r <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      Flag_AA_r <= 1'h0;
    end else begin
      if (_T_249) begin
        if (_T_251) begin
          Flag_AA_r <= 1'h1;
        end else begin
          if (_T_105) begin
            Flag_AA_r <= 1'h0;
          end
        end
      end else begin
        if (_T_260) begin
          if (_T_262) begin
            Flag_AA_r <= 1'h1;
          end else begin
            if (_T_105) begin
              Flag_AA_r <= 1'h0;
            end
          end
        end else begin
          if (_T_271) begin
            if (_T_273) begin
              Flag_AA_r <= 1'h1;
            end else begin
              if (_T_105) begin
                Flag_AA_r <= 1'h0;
              end
            end
          end else begin
            if (_T_282) begin
              if (_T_284) begin
                Flag_AA_r <= 1'h1;
              end else begin
                if (_T_105) begin
                  Flag_AA_r <= 1'h0;
                end
              end
            end else begin
              Flag_AA_r <= _GEN_53;
            end
          end
        end
      end
    end
    if (reset) begin
      Flag_AA_Valid_r <= 1'h0;
    end else begin
      if (_T_249) begin
        if (_T_251) begin
          Flag_AA_Valid_r <= 1'h1;
        end else begin
          if (_T_105) begin
            Flag_AA_Valid_r <= 1'h0;
          end
        end
      end else begin
        if (_T_260) begin
          if (_T_262) begin
            Flag_AA_Valid_r <= 1'h1;
          end else begin
            if (_T_105) begin
              Flag_AA_Valid_r <= 1'h0;
            end
          end
        end else begin
          if (_T_271) begin
            if (_T_273) begin
              Flag_AA_Valid_r <= 1'h1;
            end else begin
              if (_T_105) begin
                Flag_AA_Valid_r <= 1'h0;
              end
            end
          end else begin
            if (_T_282) begin
              Flag_AA_Valid_r <= 1'h1;
            end else begin
              if (_T_105) begin
                Flag_AA_Valid_r <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Flag_CRC_r <= 1'h0;
    end else begin
      if (_T_294) begin
        if (_T_296) begin
          Flag_CRC_r <= 1'h1;
        end else begin
          if (_T_105) begin
            Flag_CRC_r <= 1'h0;
          end
        end
      end else begin
        if (_T_305) begin
          if (_T_307) begin
            Flag_CRC_r <= 1'h1;
          end else begin
            if (_T_105) begin
              Flag_CRC_r <= 1'h0;
            end
          end
        end else begin
          if (_T_316) begin
            if (_T_318) begin
              Flag_CRC_r <= 1'h1;
            end else begin
              if (_T_105) begin
                Flag_CRC_r <= 1'h0;
              end
            end
          end else begin
            if (_T_105) begin
              Flag_CRC_r <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      Flag_CRC_Valid_r <= 1'h0;
    end else begin
      if (_T_294) begin
        if (_T_296) begin
          Flag_CRC_Valid_r <= 1'h1;
        end else begin
          if (_T_105) begin
            Flag_CRC_Valid_r <= 1'h0;
          end
        end
      end else begin
        if (_T_305) begin
          if (_T_307) begin
            Flag_CRC_Valid_r <= 1'h1;
          end else begin
            if (_T_105) begin
              Flag_CRC_Valid_r <= 1'h0;
            end
          end
        end else begin
          if (_T_316) begin
            Flag_CRC_Valid_r <= 1'h1;
          end else begin
            if (_T_105) begin
              Flag_CRC_Valid_r <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      DMA_Data_Valid_r <= 1'h0;
    end else begin
      if (_T_107) begin
        DMA_Data_Valid_r <= 1'h0;
      end else begin
        if (_T_330) begin
          DMA_Data_Valid_r <= 1'h1;
        end else begin
          if (DMA_Data_Fire_w) begin
            DMA_Data_Valid_r <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      AFIFO_Ready_r <= 1'h0;
    end else begin
      if (_T_105) begin
        AFIFO_Ready_r <= 1'h0;
      end else begin
        if (_T_106) begin
          AFIFO_Ready_r <= 1'h1;
        end else begin
          if (_T_330) begin
            AFIFO_Ready_r <= 1'h0;
          end else begin
            if (DMA_Data_Fire_w) begin
              AFIFO_Ready_r <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      data_r <= 8'h0;
    end else begin
      data_r <= _T_133;
    end
  end
endmodule
module AsyncResetRegVec_w9_i0(
  input        clock,
  input        reset,
  input  [8:0] io_d,
  output [8:0] io_q,
  input        io_en
);
  wire  reg_0_rst; // @[AsyncResetReg.scala 73:39]
  wire  reg_0_clk; // @[AsyncResetReg.scala 73:39]
  wire  reg_0_en; // @[AsyncResetReg.scala 73:39]
  wire  reg_0_q; // @[AsyncResetReg.scala 73:39]
  wire  reg_0_d; // @[AsyncResetReg.scala 73:39]
  wire  reg_1_rst; // @[AsyncResetReg.scala 73:39]
  wire  reg_1_clk; // @[AsyncResetReg.scala 73:39]
  wire  reg_1_en; // @[AsyncResetReg.scala 73:39]
  wire  reg_1_q; // @[AsyncResetReg.scala 73:39]
  wire  reg_1_d; // @[AsyncResetReg.scala 73:39]
  wire  reg_2_rst; // @[AsyncResetReg.scala 73:39]
  wire  reg_2_clk; // @[AsyncResetReg.scala 73:39]
  wire  reg_2_en; // @[AsyncResetReg.scala 73:39]
  wire  reg_2_q; // @[AsyncResetReg.scala 73:39]
  wire  reg_2_d; // @[AsyncResetReg.scala 73:39]
  wire  reg_3_rst; // @[AsyncResetReg.scala 73:39]
  wire  reg_3_clk; // @[AsyncResetReg.scala 73:39]
  wire  reg_3_en; // @[AsyncResetReg.scala 73:39]
  wire  reg_3_q; // @[AsyncResetReg.scala 73:39]
  wire  reg_3_d; // @[AsyncResetReg.scala 73:39]
  wire  reg_4_rst; // @[AsyncResetReg.scala 73:39]
  wire  reg_4_clk; // @[AsyncResetReg.scala 73:39]
  wire  reg_4_en; // @[AsyncResetReg.scala 73:39]
  wire  reg_4_q; // @[AsyncResetReg.scala 73:39]
  wire  reg_4_d; // @[AsyncResetReg.scala 73:39]
  wire  reg_5_rst; // @[AsyncResetReg.scala 73:39]
  wire  reg_5_clk; // @[AsyncResetReg.scala 73:39]
  wire  reg_5_en; // @[AsyncResetReg.scala 73:39]
  wire  reg_5_q; // @[AsyncResetReg.scala 73:39]
  wire  reg_5_d; // @[AsyncResetReg.scala 73:39]
  wire  reg_6_rst; // @[AsyncResetReg.scala 73:39]
  wire  reg_6_clk; // @[AsyncResetReg.scala 73:39]
  wire  reg_6_en; // @[AsyncResetReg.scala 73:39]
  wire  reg_6_q; // @[AsyncResetReg.scala 73:39]
  wire  reg_6_d; // @[AsyncResetReg.scala 73:39]
  wire  reg_7_rst; // @[AsyncResetReg.scala 73:39]
  wire  reg_7_clk; // @[AsyncResetReg.scala 73:39]
  wire  reg_7_en; // @[AsyncResetReg.scala 73:39]
  wire  reg_7_q; // @[AsyncResetReg.scala 73:39]
  wire  reg_7_d; // @[AsyncResetReg.scala 73:39]
  wire  reg_8_rst; // @[AsyncResetReg.scala 73:39]
  wire  reg_8_clk; // @[AsyncResetReg.scala 73:39]
  wire  reg_8_en; // @[AsyncResetReg.scala 73:39]
  wire  reg_8_q; // @[AsyncResetReg.scala 73:39]
  wire  reg_8_d; // @[AsyncResetReg.scala 73:39]
  wire  _T_5; // @[AsyncResetReg.scala 79:35]
  wire  _T_6; // @[AsyncResetReg.scala 79:35]
  wire  _T_7; // @[AsyncResetReg.scala 79:35]
  wire  _T_8; // @[AsyncResetReg.scala 79:35]
  wire  _T_9; // @[AsyncResetReg.scala 79:35]
  wire  _T_10; // @[AsyncResetReg.scala 79:35]
  wire  _T_11; // @[AsyncResetReg.scala 79:35]
  wire  _T_12; // @[AsyncResetReg.scala 79:35]
  wire  _T_13; // @[AsyncResetReg.scala 79:35]
  wire  _T_16_1; // @[AsyncResetReg.scala 85:14]
  wire  _T_16_0; // @[AsyncResetReg.scala 85:14]
  wire [1:0] _T_28; // @[AsyncResetReg.scala 85:18]
  wire  _T_16_3; // @[AsyncResetReg.scala 85:14]
  wire  _T_16_2; // @[AsyncResetReg.scala 85:14]
  wire [1:0] _T_29; // @[AsyncResetReg.scala 85:18]
  wire [3:0] _T_30; // @[AsyncResetReg.scala 85:18]
  wire  _T_16_5; // @[AsyncResetReg.scala 85:14]
  wire  _T_16_4; // @[AsyncResetReg.scala 85:14]
  wire [1:0] _T_31; // @[AsyncResetReg.scala 85:18]
  wire  _T_16_8; // @[AsyncResetReg.scala 85:14]
  wire  _T_16_7; // @[AsyncResetReg.scala 85:14]
  wire [1:0] _T_32; // @[AsyncResetReg.scala 85:18]
  wire  _T_16_6; // @[AsyncResetReg.scala 85:14]
  wire [2:0] _T_33; // @[AsyncResetReg.scala 85:18]
  wire [4:0] _T_34; // @[AsyncResetReg.scala 85:18]
  wire [8:0] _T_35; // @[AsyncResetReg.scala 85:18]
  AsyncResetReg reg_0 ( // @[AsyncResetReg.scala 73:39]
    .rst(reg_0_rst),
    .clk(reg_0_clk),
    .en(reg_0_en),
    .q(reg_0_q),
    .d(reg_0_d)
  );
  AsyncResetReg reg_1 ( // @[AsyncResetReg.scala 73:39]
    .rst(reg_1_rst),
    .clk(reg_1_clk),
    .en(reg_1_en),
    .q(reg_1_q),
    .d(reg_1_d)
  );
  AsyncResetReg reg_2 ( // @[AsyncResetReg.scala 73:39]
    .rst(reg_2_rst),
    .clk(reg_2_clk),
    .en(reg_2_en),
    .q(reg_2_q),
    .d(reg_2_d)
  );
  AsyncResetReg reg_3 ( // @[AsyncResetReg.scala 73:39]
    .rst(reg_3_rst),
    .clk(reg_3_clk),
    .en(reg_3_en),
    .q(reg_3_q),
    .d(reg_3_d)
  );
  AsyncResetReg reg_4 ( // @[AsyncResetReg.scala 73:39]
    .rst(reg_4_rst),
    .clk(reg_4_clk),
    .en(reg_4_en),
    .q(reg_4_q),
    .d(reg_4_d)
  );
  AsyncResetReg reg_5 ( // @[AsyncResetReg.scala 73:39]
    .rst(reg_5_rst),
    .clk(reg_5_clk),
    .en(reg_5_en),
    .q(reg_5_q),
    .d(reg_5_d)
  );
  AsyncResetReg reg_6 ( // @[AsyncResetReg.scala 73:39]
    .rst(reg_6_rst),
    .clk(reg_6_clk),
    .en(reg_6_en),
    .q(reg_6_q),
    .d(reg_6_d)
  );
  AsyncResetReg reg_7 ( // @[AsyncResetReg.scala 73:39]
    .rst(reg_7_rst),
    .clk(reg_7_clk),
    .en(reg_7_en),
    .q(reg_7_q),
    .d(reg_7_d)
  );
  AsyncResetReg reg_8 ( // @[AsyncResetReg.scala 73:39]
    .rst(reg_8_rst),
    .clk(reg_8_clk),
    .en(reg_8_en),
    .q(reg_8_q),
    .d(reg_8_d)
  );
  assign _T_5 = io_d[0]; // @[AsyncResetReg.scala 79:35]
  assign _T_6 = io_d[1]; // @[AsyncResetReg.scala 79:35]
  assign _T_7 = io_d[2]; // @[AsyncResetReg.scala 79:35]
  assign _T_8 = io_d[3]; // @[AsyncResetReg.scala 79:35]
  assign _T_9 = io_d[4]; // @[AsyncResetReg.scala 79:35]
  assign _T_10 = io_d[5]; // @[AsyncResetReg.scala 79:35]
  assign _T_11 = io_d[6]; // @[AsyncResetReg.scala 79:35]
  assign _T_12 = io_d[7]; // @[AsyncResetReg.scala 79:35]
  assign _T_13 = io_d[8]; // @[AsyncResetReg.scala 79:35]
  assign _T_16_1 = reg_1_q; // @[AsyncResetReg.scala 85:14]
  assign _T_16_0 = reg_0_q; // @[AsyncResetReg.scala 85:14]
  assign _T_28 = {_T_16_1,_T_16_0}; // @[AsyncResetReg.scala 85:18]
  assign _T_16_3 = reg_3_q; // @[AsyncResetReg.scala 85:14]
  assign _T_16_2 = reg_2_q; // @[AsyncResetReg.scala 85:14]
  assign _T_29 = {_T_16_3,_T_16_2}; // @[AsyncResetReg.scala 85:18]
  assign _T_30 = {_T_29,_T_28}; // @[AsyncResetReg.scala 85:18]
  assign _T_16_5 = reg_5_q; // @[AsyncResetReg.scala 85:14]
  assign _T_16_4 = reg_4_q; // @[AsyncResetReg.scala 85:14]
  assign _T_31 = {_T_16_5,_T_16_4}; // @[AsyncResetReg.scala 85:18]
  assign _T_16_8 = reg_8_q; // @[AsyncResetReg.scala 85:14]
  assign _T_16_7 = reg_7_q; // @[AsyncResetReg.scala 85:14]
  assign _T_32 = {_T_16_8,_T_16_7}; // @[AsyncResetReg.scala 85:18]
  assign _T_16_6 = reg_6_q; // @[AsyncResetReg.scala 85:14]
  assign _T_33 = {_T_32,_T_16_6}; // @[AsyncResetReg.scala 85:18]
  assign _T_34 = {_T_33,_T_31}; // @[AsyncResetReg.scala 85:18]
  assign _T_35 = {_T_34,_T_30}; // @[AsyncResetReg.scala 85:18]
  assign io_q = _T_35;
  assign reg_0_rst = reset;
  assign reg_0_clk = clock;
  assign reg_0_en = io_en;
  assign reg_0_d = _T_5;
  assign reg_1_rst = reset;
  assign reg_1_clk = clock;
  assign reg_1_en = io_en;
  assign reg_1_d = _T_6;
  assign reg_2_rst = reset;
  assign reg_2_clk = clock;
  assign reg_2_en = io_en;
  assign reg_2_d = _T_7;
  assign reg_3_rst = reset;
  assign reg_3_clk = clock;
  assign reg_3_en = io_en;
  assign reg_3_d = _T_8;
  assign reg_4_rst = reset;
  assign reg_4_clk = clock;
  assign reg_4_en = io_en;
  assign reg_4_d = _T_9;
  assign reg_5_rst = reset;
  assign reg_5_clk = clock;
  assign reg_5_en = io_en;
  assign reg_5_d = _T_10;
  assign reg_6_rst = reset;
  assign reg_6_clk = clock;
  assign reg_6_en = io_en;
  assign reg_6_d = _T_11;
  assign reg_7_rst = reset;
  assign reg_7_clk = clock;
  assign reg_7_en = io_en;
  assign reg_7_d = _T_12;
  assign reg_8_rst = reset;
  assign reg_8_clk = clock;
  assign reg_8_en = io_en;
  assign reg_8_d = _T_13;
endmodule
module AsyncResetSynchronizerShiftReg_w9_d3_i0(
  input        clock,
  input        reset,
  input  [8:0] io_d,
  output [8:0] io_q
);
  wire  sync_0_clock; // @[ShiftReg.scala 60:12]
  wire  sync_0_reset; // @[ShiftReg.scala 60:12]
  wire [8:0] sync_0_io_d; // @[ShiftReg.scala 60:12]
  wire [8:0] sync_0_io_q; // @[ShiftReg.scala 60:12]
  wire  sync_0_io_en; // @[ShiftReg.scala 60:12]
  wire  sync_1_clock; // @[ShiftReg.scala 60:12]
  wire  sync_1_reset; // @[ShiftReg.scala 60:12]
  wire [8:0] sync_1_io_d; // @[ShiftReg.scala 60:12]
  wire [8:0] sync_1_io_q; // @[ShiftReg.scala 60:12]
  wire  sync_1_io_en; // @[ShiftReg.scala 60:12]
  wire  sync_2_clock; // @[ShiftReg.scala 60:12]
  wire  sync_2_reset; // @[ShiftReg.scala 60:12]
  wire [8:0] sync_2_io_d; // @[ShiftReg.scala 60:12]
  wire [8:0] sync_2_io_q; // @[ShiftReg.scala 60:12]
  wire  sync_2_io_en; // @[ShiftReg.scala 60:12]
  AsyncResetRegVec_w9_i0 sync_0 ( // @[ShiftReg.scala 60:12]
    .clock(sync_0_clock),
    .reset(sync_0_reset),
    .io_d(sync_0_io_d),
    .io_q(sync_0_io_q),
    .io_en(sync_0_io_en)
  );
  AsyncResetRegVec_w9_i0 sync_1 ( // @[ShiftReg.scala 60:12]
    .clock(sync_1_clock),
    .reset(sync_1_reset),
    .io_d(sync_1_io_d),
    .io_q(sync_1_io_q),
    .io_en(sync_1_io_en)
  );
  AsyncResetRegVec_w9_i0 sync_2 ( // @[ShiftReg.scala 60:12]
    .clock(sync_2_clock),
    .reset(sync_2_reset),
    .io_d(sync_2_io_d),
    .io_q(sync_2_io_q),
    .io_en(sync_2_io_en)
  );
  assign io_q = sync_0_io_q;
  assign sync_0_clock = clock;
  assign sync_0_reset = reset;
  assign sync_0_io_d = sync_1_io_q;
  assign sync_0_io_en = 1'h1;
  assign sync_1_clock = clock;
  assign sync_1_reset = reset;
  assign sync_1_io_d = sync_2_io_q;
  assign sync_1_io_en = 1'h1;
  assign sync_2_clock = clock;
  assign sync_2_reset = reset;
  assign sync_2_io_d = io_d;
  assign sync_2_io_en = 1'h1;
endmodule
module AsyncResetRegVec_w1_i0(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q,
  input   io_en
);
  wire  reg_0_rst; // @[AsyncResetReg.scala 73:39]
  wire  reg_0_clk; // @[AsyncResetReg.scala 73:39]
  wire  reg_0_en; // @[AsyncResetReg.scala 73:39]
  wire  reg_0_q; // @[AsyncResetReg.scala 73:39]
  wire  reg_0_d; // @[AsyncResetReg.scala 73:39]
  wire  _T_8_0; // @[AsyncResetReg.scala 85:14]
  AsyncResetReg reg_0 ( // @[AsyncResetReg.scala 73:39]
    .rst(reg_0_rst),
    .clk(reg_0_clk),
    .en(reg_0_en),
    .q(reg_0_q),
    .d(reg_0_d)
  );
  assign _T_8_0 = reg_0_q; // @[AsyncResetReg.scala 85:14]
  assign io_q = _T_8_0;
  assign reg_0_rst = reset;
  assign reg_0_clk = clock;
  assign reg_0_en = io_en;
  assign reg_0_d = io_d;
endmodule
module AsyncResetSynchronizerShiftReg_w1_d4_i0(
  input   clock,
  input   reset,
  output  io_q
);
  wire  sync_0_clock; // @[ShiftReg.scala 60:12]
  wire  sync_0_reset; // @[ShiftReg.scala 60:12]
  wire  sync_0_io_d; // @[ShiftReg.scala 60:12]
  wire  sync_0_io_q; // @[ShiftReg.scala 60:12]
  wire  sync_0_io_en; // @[ShiftReg.scala 60:12]
  wire  sync_1_clock; // @[ShiftReg.scala 60:12]
  wire  sync_1_reset; // @[ShiftReg.scala 60:12]
  wire  sync_1_io_d; // @[ShiftReg.scala 60:12]
  wire  sync_1_io_q; // @[ShiftReg.scala 60:12]
  wire  sync_1_io_en; // @[ShiftReg.scala 60:12]
  wire  sync_2_clock; // @[ShiftReg.scala 60:12]
  wire  sync_2_reset; // @[ShiftReg.scala 60:12]
  wire  sync_2_io_d; // @[ShiftReg.scala 60:12]
  wire  sync_2_io_q; // @[ShiftReg.scala 60:12]
  wire  sync_2_io_en; // @[ShiftReg.scala 60:12]
  wire  sync_3_clock; // @[ShiftReg.scala 60:12]
  wire  sync_3_reset; // @[ShiftReg.scala 60:12]
  wire  sync_3_io_d; // @[ShiftReg.scala 60:12]
  wire  sync_3_io_q; // @[ShiftReg.scala 60:12]
  wire  sync_3_io_en; // @[ShiftReg.scala 60:12]
  AsyncResetRegVec_w1_i0 sync_0 ( // @[ShiftReg.scala 60:12]
    .clock(sync_0_clock),
    .reset(sync_0_reset),
    .io_d(sync_0_io_d),
    .io_q(sync_0_io_q),
    .io_en(sync_0_io_en)
  );
  AsyncResetRegVec_w1_i0 sync_1 ( // @[ShiftReg.scala 60:12]
    .clock(sync_1_clock),
    .reset(sync_1_reset),
    .io_d(sync_1_io_d),
    .io_q(sync_1_io_q),
    .io_en(sync_1_io_en)
  );
  AsyncResetRegVec_w1_i0 sync_2 ( // @[ShiftReg.scala 60:12]
    .clock(sync_2_clock),
    .reset(sync_2_reset),
    .io_d(sync_2_io_d),
    .io_q(sync_2_io_q),
    .io_en(sync_2_io_en)
  );
  AsyncResetRegVec_w1_i0 sync_3 ( // @[ShiftReg.scala 60:12]
    .clock(sync_3_clock),
    .reset(sync_3_reset),
    .io_d(sync_3_io_d),
    .io_q(sync_3_io_q),
    .io_en(sync_3_io_en)
  );
  assign io_q = sync_0_io_q;
  assign sync_0_clock = clock;
  assign sync_0_reset = reset;
  assign sync_0_io_d = sync_1_io_q;
  assign sync_0_io_en = 1'h1;
  assign sync_1_clock = clock;
  assign sync_1_reset = reset;
  assign sync_1_io_d = sync_2_io_q;
  assign sync_1_io_en = 1'h1;
  assign sync_2_clock = clock;
  assign sync_2_reset = reset;
  assign sync_2_io_d = sync_3_io_q;
  assign sync_2_io_en = 1'h1;
  assign sync_3_clock = clock;
  assign sync_3_reset = reset;
  assign sync_3_io_d = 1'h1;
  assign sync_3_io_en = 1'h1;
endmodule
module AsyncValidSync(
  input   clock,
  input   reset,
  output  io_out
);
  wire  source_valid_clock; // @[ShiftReg.scala 47:23]
  wire  source_valid_reset; // @[ShiftReg.scala 47:23]
  wire  source_valid_io_q; // @[ShiftReg.scala 47:23]
  wire  _T_5; // @[ShiftReg.scala 50:24]
  AsyncResetSynchronizerShiftReg_w1_d4_i0 source_valid ( // @[ShiftReg.scala 47:23]
    .clock(source_valid_clock),
    .reset(source_valid_reset),
    .io_q(source_valid_io_q)
  );
  assign _T_5 = source_valid_io_q; // @[ShiftReg.scala 50:24]
  assign io_out = _T_5;
  assign source_valid_clock = clock;
  assign source_valid_reset = reset;
endmodule
module AsyncResetSynchronizerShiftReg_w1_d1_i0(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q
);
  wire  sync_0_clock; // @[ShiftReg.scala 60:12]
  wire  sync_0_reset; // @[ShiftReg.scala 60:12]
  wire  sync_0_io_d; // @[ShiftReg.scala 60:12]
  wire  sync_0_io_q; // @[ShiftReg.scala 60:12]
  wire  sync_0_io_en; // @[ShiftReg.scala 60:12]
  AsyncResetRegVec_w1_i0 sync_0 ( // @[ShiftReg.scala 60:12]
    .clock(sync_0_clock),
    .reset(sync_0_reset),
    .io_d(sync_0_io_d),
    .io_q(sync_0_io_q),
    .io_en(sync_0_io_en)
  );
  assign io_q = sync_0_io_q;
  assign sync_0_clock = clock;
  assign sync_0_reset = reset;
  assign sync_0_io_d = io_d;
  assign sync_0_io_en = 1'h1;
endmodule
module AsyncValidSync_1(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  sink_extend_clock; // @[ShiftReg.scala 47:23]
  wire  sink_extend_reset; // @[ShiftReg.scala 47:23]
  wire  sink_extend_io_d; // @[ShiftReg.scala 47:23]
  wire  sink_extend_io_q; // @[ShiftReg.scala 47:23]
  wire  _T_5; // @[ShiftReg.scala 50:24]
  AsyncResetSynchronizerShiftReg_w1_d1_i0 sink_extend ( // @[ShiftReg.scala 47:23]
    .clock(sink_extend_clock),
    .reset(sink_extend_reset),
    .io_d(sink_extend_io_d),
    .io_q(sink_extend_io_q)
  );
  assign _T_5 = sink_extend_io_q; // @[ShiftReg.scala 50:24]
  assign io_out = _T_5;
  assign sink_extend_clock = clock;
  assign sink_extend_reset = reset;
  assign sink_extend_io_d = io_in;
endmodule
module AsyncResetSynchronizerShiftReg_w1_d3_i0(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q
);
  wire  sync_0_clock; // @[ShiftReg.scala 60:12]
  wire  sync_0_reset; // @[ShiftReg.scala 60:12]
  wire  sync_0_io_d; // @[ShiftReg.scala 60:12]
  wire  sync_0_io_q; // @[ShiftReg.scala 60:12]
  wire  sync_0_io_en; // @[ShiftReg.scala 60:12]
  wire  sync_1_clock; // @[ShiftReg.scala 60:12]
  wire  sync_1_reset; // @[ShiftReg.scala 60:12]
  wire  sync_1_io_d; // @[ShiftReg.scala 60:12]
  wire  sync_1_io_q; // @[ShiftReg.scala 60:12]
  wire  sync_1_io_en; // @[ShiftReg.scala 60:12]
  wire  sync_2_clock; // @[ShiftReg.scala 60:12]
  wire  sync_2_reset; // @[ShiftReg.scala 60:12]
  wire  sync_2_io_d; // @[ShiftReg.scala 60:12]
  wire  sync_2_io_q; // @[ShiftReg.scala 60:12]
  wire  sync_2_io_en; // @[ShiftReg.scala 60:12]
  AsyncResetRegVec_w1_i0 sync_0 ( // @[ShiftReg.scala 60:12]
    .clock(sync_0_clock),
    .reset(sync_0_reset),
    .io_d(sync_0_io_d),
    .io_q(sync_0_io_q),
    .io_en(sync_0_io_en)
  );
  AsyncResetRegVec_w1_i0 sync_1 ( // @[ShiftReg.scala 60:12]
    .clock(sync_1_clock),
    .reset(sync_1_reset),
    .io_d(sync_1_io_d),
    .io_q(sync_1_io_q),
    .io_en(sync_1_io_en)
  );
  AsyncResetRegVec_w1_i0 sync_2 ( // @[ShiftReg.scala 60:12]
    .clock(sync_2_clock),
    .reset(sync_2_reset),
    .io_d(sync_2_io_d),
    .io_q(sync_2_io_q),
    .io_en(sync_2_io_en)
  );
  assign io_q = sync_0_io_q;
  assign sync_0_clock = clock;
  assign sync_0_reset = reset;
  assign sync_0_io_d = sync_1_io_q;
  assign sync_0_io_en = 1'h1;
  assign sync_1_clock = clock;
  assign sync_1_reset = reset;
  assign sync_1_io_d = sync_2_io_q;
  assign sync_1_io_en = 1'h1;
  assign sync_2_clock = clock;
  assign sync_2_reset = reset;
  assign sync_2_io_d = io_d;
  assign sync_2_io_en = 1'h1;
endmodule
module AsyncValidSync_2(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  sink_valid_clock; // @[ShiftReg.scala 47:23]
  wire  sink_valid_reset; // @[ShiftReg.scala 47:23]
  wire  sink_valid_io_d; // @[ShiftReg.scala 47:23]
  wire  sink_valid_io_q; // @[ShiftReg.scala 47:23]
  wire  _T_5; // @[ShiftReg.scala 50:24]
  AsyncResetSynchronizerShiftReg_w1_d3_i0 sink_valid ( // @[ShiftReg.scala 47:23]
    .clock(sink_valid_clock),
    .reset(sink_valid_reset),
    .io_d(sink_valid_io_d),
    .io_q(sink_valid_io_q)
  );
  assign _T_5 = sink_valid_io_q; // @[ShiftReg.scala 50:24]
  assign io_out = _T_5;
  assign sink_valid_clock = clock;
  assign sink_valid_reset = reset;
  assign sink_valid_io_d = io_in;
endmodule
module AsyncQueueSource(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input        io_enq_bits,
  input  [8:0] io_ridx,
  output [8:0] io_widx,
  output       io_mem_0,
  output       io_mem_1,
  output       io_mem_2,
  output       io_mem_3,
  output       io_mem_4,
  output       io_mem_5,
  output       io_mem_6,
  output       io_mem_7,
  output       io_mem_8,
  output       io_mem_9,
  output       io_mem_10,
  output       io_mem_11,
  output       io_mem_12,
  output       io_mem_13,
  output       io_mem_14,
  output       io_mem_15,
  output       io_mem_16,
  output       io_mem_17,
  output       io_mem_18,
  output       io_mem_19,
  output       io_mem_20,
  output       io_mem_21,
  output       io_mem_22,
  output       io_mem_23,
  output       io_mem_24,
  output       io_mem_25,
  output       io_mem_26,
  output       io_mem_27,
  output       io_mem_28,
  output       io_mem_29,
  output       io_mem_30,
  output       io_mem_31,
  output       io_mem_32,
  output       io_mem_33,
  output       io_mem_34,
  output       io_mem_35,
  output       io_mem_36,
  output       io_mem_37,
  output       io_mem_38,
  output       io_mem_39,
  output       io_mem_40,
  output       io_mem_41,
  output       io_mem_42,
  output       io_mem_43,
  output       io_mem_44,
  output       io_mem_45,
  output       io_mem_46,
  output       io_mem_47,
  output       io_mem_48,
  output       io_mem_49,
  output       io_mem_50,
  output       io_mem_51,
  output       io_mem_52,
  output       io_mem_53,
  output       io_mem_54,
  output       io_mem_55,
  output       io_mem_56,
  output       io_mem_57,
  output       io_mem_58,
  output       io_mem_59,
  output       io_mem_60,
  output       io_mem_61,
  output       io_mem_62,
  output       io_mem_63,
  output       io_mem_64,
  output       io_mem_65,
  output       io_mem_66,
  output       io_mem_67,
  output       io_mem_68,
  output       io_mem_69,
  output       io_mem_70,
  output       io_mem_71,
  output       io_mem_72,
  output       io_mem_73,
  output       io_mem_74,
  output       io_mem_75,
  output       io_mem_76,
  output       io_mem_77,
  output       io_mem_78,
  output       io_mem_79,
  output       io_mem_80,
  output       io_mem_81,
  output       io_mem_82,
  output       io_mem_83,
  output       io_mem_84,
  output       io_mem_85,
  output       io_mem_86,
  output       io_mem_87,
  output       io_mem_88,
  output       io_mem_89,
  output       io_mem_90,
  output       io_mem_91,
  output       io_mem_92,
  output       io_mem_93,
  output       io_mem_94,
  output       io_mem_95,
  output       io_mem_96,
  output       io_mem_97,
  output       io_mem_98,
  output       io_mem_99,
  output       io_mem_100,
  output       io_mem_101,
  output       io_mem_102,
  output       io_mem_103,
  output       io_mem_104,
  output       io_mem_105,
  output       io_mem_106,
  output       io_mem_107,
  output       io_mem_108,
  output       io_mem_109,
  output       io_mem_110,
  output       io_mem_111,
  output       io_mem_112,
  output       io_mem_113,
  output       io_mem_114,
  output       io_mem_115,
  output       io_mem_116,
  output       io_mem_117,
  output       io_mem_118,
  output       io_mem_119,
  output       io_mem_120,
  output       io_mem_121,
  output       io_mem_122,
  output       io_mem_123,
  output       io_mem_124,
  output       io_mem_125,
  output       io_mem_126,
  output       io_mem_127,
  output       io_mem_128,
  output       io_mem_129,
  output       io_mem_130,
  output       io_mem_131,
  output       io_mem_132,
  output       io_mem_133,
  output       io_mem_134,
  output       io_mem_135,
  output       io_mem_136,
  output       io_mem_137,
  output       io_mem_138,
  output       io_mem_139,
  output       io_mem_140,
  output       io_mem_141,
  output       io_mem_142,
  output       io_mem_143,
  output       io_mem_144,
  output       io_mem_145,
  output       io_mem_146,
  output       io_mem_147,
  output       io_mem_148,
  output       io_mem_149,
  output       io_mem_150,
  output       io_mem_151,
  output       io_mem_152,
  output       io_mem_153,
  output       io_mem_154,
  output       io_mem_155,
  output       io_mem_156,
  output       io_mem_157,
  output       io_mem_158,
  output       io_mem_159,
  output       io_mem_160,
  output       io_mem_161,
  output       io_mem_162,
  output       io_mem_163,
  output       io_mem_164,
  output       io_mem_165,
  output       io_mem_166,
  output       io_mem_167,
  output       io_mem_168,
  output       io_mem_169,
  output       io_mem_170,
  output       io_mem_171,
  output       io_mem_172,
  output       io_mem_173,
  output       io_mem_174,
  output       io_mem_175,
  output       io_mem_176,
  output       io_mem_177,
  output       io_mem_178,
  output       io_mem_179,
  output       io_mem_180,
  output       io_mem_181,
  output       io_mem_182,
  output       io_mem_183,
  output       io_mem_184,
  output       io_mem_185,
  output       io_mem_186,
  output       io_mem_187,
  output       io_mem_188,
  output       io_mem_189,
  output       io_mem_190,
  output       io_mem_191,
  output       io_mem_192,
  output       io_mem_193,
  output       io_mem_194,
  output       io_mem_195,
  output       io_mem_196,
  output       io_mem_197,
  output       io_mem_198,
  output       io_mem_199,
  output       io_mem_200,
  output       io_mem_201,
  output       io_mem_202,
  output       io_mem_203,
  output       io_mem_204,
  output       io_mem_205,
  output       io_mem_206,
  output       io_mem_207,
  output       io_mem_208,
  output       io_mem_209,
  output       io_mem_210,
  output       io_mem_211,
  output       io_mem_212,
  output       io_mem_213,
  output       io_mem_214,
  output       io_mem_215,
  output       io_mem_216,
  output       io_mem_217,
  output       io_mem_218,
  output       io_mem_219,
  output       io_mem_220,
  output       io_mem_221,
  output       io_mem_222,
  output       io_mem_223,
  output       io_mem_224,
  output       io_mem_225,
  output       io_mem_226,
  output       io_mem_227,
  output       io_mem_228,
  output       io_mem_229,
  output       io_mem_230,
  output       io_mem_231,
  output       io_mem_232,
  output       io_mem_233,
  output       io_mem_234,
  output       io_mem_235,
  output       io_mem_236,
  output       io_mem_237,
  output       io_mem_238,
  output       io_mem_239,
  output       io_mem_240,
  output       io_mem_241,
  output       io_mem_242,
  output       io_mem_243,
  output       io_mem_244,
  output       io_mem_245,
  output       io_mem_246,
  output       io_mem_247,
  output       io_mem_248,
  output       io_mem_249,
  output       io_mem_250,
  output       io_mem_251,
  output       io_mem_252,
  output       io_mem_253,
  output       io_mem_254,
  output       io_mem_255,
  input        io_sink_reset_n,
  input        io_ridx_valid,
  output       io_widx_valid
);
  reg  mem_0; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_0;
  reg  mem_1; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_1;
  reg  mem_2; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_2;
  reg  mem_3; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_3;
  reg  mem_4; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_4;
  reg  mem_5; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_5;
  reg  mem_6; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_6;
  reg  mem_7; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_7;
  reg  mem_8; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_8;
  reg  mem_9; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_9;
  reg  mem_10; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_10;
  reg  mem_11; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_11;
  reg  mem_12; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_12;
  reg  mem_13; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_13;
  reg  mem_14; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_14;
  reg  mem_15; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_15;
  reg  mem_16; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_16;
  reg  mem_17; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_17;
  reg  mem_18; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_18;
  reg  mem_19; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_19;
  reg  mem_20; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_20;
  reg  mem_21; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_21;
  reg  mem_22; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_22;
  reg  mem_23; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_23;
  reg  mem_24; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_24;
  reg  mem_25; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_25;
  reg  mem_26; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_26;
  reg  mem_27; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_27;
  reg  mem_28; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_28;
  reg  mem_29; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_29;
  reg  mem_30; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_30;
  reg  mem_31; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_31;
  reg  mem_32; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_32;
  reg  mem_33; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_33;
  reg  mem_34; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_34;
  reg  mem_35; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_35;
  reg  mem_36; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_36;
  reg  mem_37; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_37;
  reg  mem_38; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_38;
  reg  mem_39; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_39;
  reg  mem_40; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_40;
  reg  mem_41; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_41;
  reg  mem_42; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_42;
  reg  mem_43; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_43;
  reg  mem_44; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_44;
  reg  mem_45; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_45;
  reg  mem_46; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_46;
  reg  mem_47; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_47;
  reg  mem_48; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_48;
  reg  mem_49; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_49;
  reg  mem_50; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_50;
  reg  mem_51; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_51;
  reg  mem_52; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_52;
  reg  mem_53; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_53;
  reg  mem_54; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_54;
  reg  mem_55; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_55;
  reg  mem_56; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_56;
  reg  mem_57; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_57;
  reg  mem_58; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_58;
  reg  mem_59; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_59;
  reg  mem_60; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_60;
  reg  mem_61; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_61;
  reg  mem_62; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_62;
  reg  mem_63; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_63;
  reg  mem_64; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_64;
  reg  mem_65; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_65;
  reg  mem_66; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_66;
  reg  mem_67; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_67;
  reg  mem_68; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_68;
  reg  mem_69; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_69;
  reg  mem_70; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_70;
  reg  mem_71; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_71;
  reg  mem_72; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_72;
  reg  mem_73; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_73;
  reg  mem_74; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_74;
  reg  mem_75; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_75;
  reg  mem_76; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_76;
  reg  mem_77; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_77;
  reg  mem_78; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_78;
  reg  mem_79; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_79;
  reg  mem_80; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_80;
  reg  mem_81; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_81;
  reg  mem_82; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_82;
  reg  mem_83; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_83;
  reg  mem_84; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_84;
  reg  mem_85; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_85;
  reg  mem_86; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_86;
  reg  mem_87; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_87;
  reg  mem_88; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_88;
  reg  mem_89; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_89;
  reg  mem_90; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_90;
  reg  mem_91; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_91;
  reg  mem_92; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_92;
  reg  mem_93; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_93;
  reg  mem_94; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_94;
  reg  mem_95; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_95;
  reg  mem_96; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_96;
  reg  mem_97; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_97;
  reg  mem_98; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_98;
  reg  mem_99; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_99;
  reg  mem_100; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_100;
  reg  mem_101; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_101;
  reg  mem_102; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_102;
  reg  mem_103; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_103;
  reg  mem_104; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_104;
  reg  mem_105; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_105;
  reg  mem_106; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_106;
  reg  mem_107; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_107;
  reg  mem_108; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_108;
  reg  mem_109; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_109;
  reg  mem_110; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_110;
  reg  mem_111; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_111;
  reg  mem_112; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_112;
  reg  mem_113; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_113;
  reg  mem_114; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_114;
  reg  mem_115; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_115;
  reg  mem_116; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_116;
  reg  mem_117; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_117;
  reg  mem_118; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_118;
  reg  mem_119; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_119;
  reg  mem_120; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_120;
  reg  mem_121; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_121;
  reg  mem_122; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_122;
  reg  mem_123; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_123;
  reg  mem_124; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_124;
  reg  mem_125; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_125;
  reg  mem_126; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_126;
  reg  mem_127; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_127;
  reg  mem_128; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_128;
  reg  mem_129; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_129;
  reg  mem_130; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_130;
  reg  mem_131; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_131;
  reg  mem_132; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_132;
  reg  mem_133; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_133;
  reg  mem_134; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_134;
  reg  mem_135; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_135;
  reg  mem_136; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_136;
  reg  mem_137; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_137;
  reg  mem_138; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_138;
  reg  mem_139; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_139;
  reg  mem_140; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_140;
  reg  mem_141; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_141;
  reg  mem_142; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_142;
  reg  mem_143; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_143;
  reg  mem_144; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_144;
  reg  mem_145; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_145;
  reg  mem_146; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_146;
  reg  mem_147; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_147;
  reg  mem_148; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_148;
  reg  mem_149; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_149;
  reg  mem_150; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_150;
  reg  mem_151; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_151;
  reg  mem_152; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_152;
  reg  mem_153; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_153;
  reg  mem_154; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_154;
  reg  mem_155; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_155;
  reg  mem_156; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_156;
  reg  mem_157; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_157;
  reg  mem_158; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_158;
  reg  mem_159; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_159;
  reg  mem_160; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_160;
  reg  mem_161; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_161;
  reg  mem_162; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_162;
  reg  mem_163; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_163;
  reg  mem_164; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_164;
  reg  mem_165; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_165;
  reg  mem_166; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_166;
  reg  mem_167; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_167;
  reg  mem_168; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_168;
  reg  mem_169; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_169;
  reg  mem_170; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_170;
  reg  mem_171; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_171;
  reg  mem_172; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_172;
  reg  mem_173; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_173;
  reg  mem_174; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_174;
  reg  mem_175; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_175;
  reg  mem_176; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_176;
  reg  mem_177; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_177;
  reg  mem_178; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_178;
  reg  mem_179; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_179;
  reg  mem_180; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_180;
  reg  mem_181; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_181;
  reg  mem_182; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_182;
  reg  mem_183; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_183;
  reg  mem_184; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_184;
  reg  mem_185; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_185;
  reg  mem_186; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_186;
  reg  mem_187; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_187;
  reg  mem_188; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_188;
  reg  mem_189; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_189;
  reg  mem_190; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_190;
  reg  mem_191; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_191;
  reg  mem_192; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_192;
  reg  mem_193; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_193;
  reg  mem_194; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_194;
  reg  mem_195; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_195;
  reg  mem_196; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_196;
  reg  mem_197; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_197;
  reg  mem_198; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_198;
  reg  mem_199; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_199;
  reg  mem_200; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_200;
  reg  mem_201; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_201;
  reg  mem_202; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_202;
  reg  mem_203; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_203;
  reg  mem_204; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_204;
  reg  mem_205; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_205;
  reg  mem_206; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_206;
  reg  mem_207; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_207;
  reg  mem_208; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_208;
  reg  mem_209; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_209;
  reg  mem_210; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_210;
  reg  mem_211; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_211;
  reg  mem_212; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_212;
  reg  mem_213; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_213;
  reg  mem_214; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_214;
  reg  mem_215; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_215;
  reg  mem_216; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_216;
  reg  mem_217; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_217;
  reg  mem_218; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_218;
  reg  mem_219; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_219;
  reg  mem_220; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_220;
  reg  mem_221; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_221;
  reg  mem_222; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_222;
  reg  mem_223; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_223;
  reg  mem_224; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_224;
  reg  mem_225; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_225;
  reg  mem_226; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_226;
  reg  mem_227; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_227;
  reg  mem_228; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_228;
  reg  mem_229; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_229;
  reg  mem_230; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_230;
  reg  mem_231; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_231;
  reg  mem_232; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_232;
  reg  mem_233; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_233;
  reg  mem_234; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_234;
  reg  mem_235; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_235;
  reg  mem_236; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_236;
  reg  mem_237; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_237;
  reg  mem_238; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_238;
  reg  mem_239; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_239;
  reg  mem_240; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_240;
  reg  mem_241; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_241;
  reg  mem_242; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_242;
  reg  mem_243; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_243;
  reg  mem_244; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_244;
  reg  mem_245; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_245;
  reg  mem_246; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_246;
  reg  mem_247; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_247;
  reg  mem_248; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_248;
  reg  mem_249; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_249;
  reg  mem_250; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_250;
  reg  mem_251; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_251;
  reg  mem_252; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_252;
  reg  mem_253; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_253;
  reg  mem_254; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_254;
  reg  mem_255; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_255;
  wire  widx_bin_clock; // @[AsyncResetReg.scala 110:21]
  wire  widx_bin_reset; // @[AsyncResetReg.scala 110:21]
  wire [8:0] widx_bin_io_d; // @[AsyncResetReg.scala 110:21]
  wire [8:0] widx_bin_io_q; // @[AsyncResetReg.scala 110:21]
  wire  widx_bin_io_en; // @[AsyncResetReg.scala 110:21]
  wire  ridx_gray_clock; // @[ShiftReg.scala 47:23]
  wire  ridx_gray_reset; // @[ShiftReg.scala 47:23]
  wire [8:0] ridx_gray_io_d; // @[ShiftReg.scala 47:23]
  wire [8:0] ridx_gray_io_q; // @[ShiftReg.scala 47:23]
  wire  ready_reg_clock; // @[AsyncResetReg.scala 110:21]
  wire  ready_reg_reset; // @[AsyncResetReg.scala 110:21]
  wire  ready_reg_io_d; // @[AsyncResetReg.scala 110:21]
  wire  ready_reg_io_q; // @[AsyncResetReg.scala 110:21]
  wire  ready_reg_io_en; // @[AsyncResetReg.scala 110:21]
  wire  widx_gray_clock; // @[AsyncResetReg.scala 110:21]
  wire  widx_gray_reset; // @[AsyncResetReg.scala 110:21]
  wire [8:0] widx_gray_io_d; // @[AsyncResetReg.scala 110:21]
  wire [8:0] widx_gray_io_q; // @[AsyncResetReg.scala 110:21]
  wire  widx_gray_io_en; // @[AsyncResetReg.scala 110:21]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 59:30]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 59:30]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 59:30]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 60:30]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 60:30]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 60:30]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 60:30]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 61:30]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 61:30]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 61:30]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 61:30]
  wire  _T_536; // @[Decoupled.scala 30:37]
  wire  sink_ready;
  wire  _T_538; // @[AsyncQueue.scala 42:49]
  wire [8:0] _GEN_513; // @[AsyncQueue.scala 11:47]
  wire [9:0] _T_543; // @[AsyncQueue.scala 11:47]
  wire [8:0] _T_544; // @[AsyncQueue.scala 11:47]
  wire [8:0] _T_545; // @[AsyncQueue.scala 11:23]
  wire [8:0] _T_547; // @[AsyncQueue.scala 12:32]
  wire [8:0] widx; // @[AsyncQueue.scala 12:17]
  wire [8:0] ridx; // @[ShiftReg.scala 50:24]
  wire [8:0] _T_550; // @[AsyncQueue.scala 44:44]
  wire  _T_551; // @[AsyncQueue.scala 44:34]
  wire  ready; // @[AsyncQueue.scala 44:26]
  wire [7:0] _T_552; // @[AsyncQueue.scala 46:51]
  wire  _T_553; // @[AsyncQueue.scala 46:73]
  wire [7:0] _GEN_514; // @[AsyncQueue.scala 46:86]
  wire [7:0] _T_554; // @[AsyncQueue.scala 46:86]
  wire [7:0] index; // @[AsyncQueue.scala 46:63]
  wire  _GEN_1; // @[AsyncQueue.scala 47:37]
  wire  _GEN_2; // @[AsyncQueue.scala 47:37]
  wire  _GEN_3; // @[AsyncQueue.scala 47:37]
  wire  _GEN_4; // @[AsyncQueue.scala 47:37]
  wire  _GEN_5; // @[AsyncQueue.scala 47:37]
  wire  _GEN_6; // @[AsyncQueue.scala 47:37]
  wire  _GEN_7; // @[AsyncQueue.scala 47:37]
  wire  _GEN_8; // @[AsyncQueue.scala 47:37]
  wire  _GEN_9; // @[AsyncQueue.scala 47:37]
  wire  _GEN_10; // @[AsyncQueue.scala 47:37]
  wire  _GEN_11; // @[AsyncQueue.scala 47:37]
  wire  _GEN_12; // @[AsyncQueue.scala 47:37]
  wire  _GEN_13; // @[AsyncQueue.scala 47:37]
  wire  _GEN_14; // @[AsyncQueue.scala 47:37]
  wire  _GEN_15; // @[AsyncQueue.scala 47:37]
  wire  _GEN_16; // @[AsyncQueue.scala 47:37]
  wire  _GEN_17; // @[AsyncQueue.scala 47:37]
  wire  _GEN_18; // @[AsyncQueue.scala 47:37]
  wire  _GEN_19; // @[AsyncQueue.scala 47:37]
  wire  _GEN_20; // @[AsyncQueue.scala 47:37]
  wire  _GEN_21; // @[AsyncQueue.scala 47:37]
  wire  _GEN_22; // @[AsyncQueue.scala 47:37]
  wire  _GEN_23; // @[AsyncQueue.scala 47:37]
  wire  _GEN_24; // @[AsyncQueue.scala 47:37]
  wire  _GEN_25; // @[AsyncQueue.scala 47:37]
  wire  _GEN_26; // @[AsyncQueue.scala 47:37]
  wire  _GEN_27; // @[AsyncQueue.scala 47:37]
  wire  _GEN_28; // @[AsyncQueue.scala 47:37]
  wire  _GEN_29; // @[AsyncQueue.scala 47:37]
  wire  _GEN_30; // @[AsyncQueue.scala 47:37]
  wire  _GEN_31; // @[AsyncQueue.scala 47:37]
  wire  _GEN_32; // @[AsyncQueue.scala 47:37]
  wire  _GEN_33; // @[AsyncQueue.scala 47:37]
  wire  _GEN_34; // @[AsyncQueue.scala 47:37]
  wire  _GEN_35; // @[AsyncQueue.scala 47:37]
  wire  _GEN_36; // @[AsyncQueue.scala 47:37]
  wire  _GEN_37; // @[AsyncQueue.scala 47:37]
  wire  _GEN_38; // @[AsyncQueue.scala 47:37]
  wire  _GEN_39; // @[AsyncQueue.scala 47:37]
  wire  _GEN_40; // @[AsyncQueue.scala 47:37]
  wire  _GEN_41; // @[AsyncQueue.scala 47:37]
  wire  _GEN_42; // @[AsyncQueue.scala 47:37]
  wire  _GEN_43; // @[AsyncQueue.scala 47:37]
  wire  _GEN_44; // @[AsyncQueue.scala 47:37]
  wire  _GEN_45; // @[AsyncQueue.scala 47:37]
  wire  _GEN_46; // @[AsyncQueue.scala 47:37]
  wire  _GEN_47; // @[AsyncQueue.scala 47:37]
  wire  _GEN_48; // @[AsyncQueue.scala 47:37]
  wire  _GEN_49; // @[AsyncQueue.scala 47:37]
  wire  _GEN_50; // @[AsyncQueue.scala 47:37]
  wire  _GEN_51; // @[AsyncQueue.scala 47:37]
  wire  _GEN_52; // @[AsyncQueue.scala 47:37]
  wire  _GEN_53; // @[AsyncQueue.scala 47:37]
  wire  _GEN_54; // @[AsyncQueue.scala 47:37]
  wire  _GEN_55; // @[AsyncQueue.scala 47:37]
  wire  _GEN_56; // @[AsyncQueue.scala 47:37]
  wire  _GEN_57; // @[AsyncQueue.scala 47:37]
  wire  _GEN_58; // @[AsyncQueue.scala 47:37]
  wire  _GEN_59; // @[AsyncQueue.scala 47:37]
  wire  _GEN_60; // @[AsyncQueue.scala 47:37]
  wire  _GEN_61; // @[AsyncQueue.scala 47:37]
  wire  _GEN_62; // @[AsyncQueue.scala 47:37]
  wire  _GEN_63; // @[AsyncQueue.scala 47:37]
  wire  _GEN_64; // @[AsyncQueue.scala 47:37]
  wire  _GEN_65; // @[AsyncQueue.scala 47:37]
  wire  _GEN_66; // @[AsyncQueue.scala 47:37]
  wire  _GEN_67; // @[AsyncQueue.scala 47:37]
  wire  _GEN_68; // @[AsyncQueue.scala 47:37]
  wire  _GEN_69; // @[AsyncQueue.scala 47:37]
  wire  _GEN_70; // @[AsyncQueue.scala 47:37]
  wire  _GEN_71; // @[AsyncQueue.scala 47:37]
  wire  _GEN_72; // @[AsyncQueue.scala 47:37]
  wire  _GEN_73; // @[AsyncQueue.scala 47:37]
  wire  _GEN_74; // @[AsyncQueue.scala 47:37]
  wire  _GEN_75; // @[AsyncQueue.scala 47:37]
  wire  _GEN_76; // @[AsyncQueue.scala 47:37]
  wire  _GEN_77; // @[AsyncQueue.scala 47:37]
  wire  _GEN_78; // @[AsyncQueue.scala 47:37]
  wire  _GEN_79; // @[AsyncQueue.scala 47:37]
  wire  _GEN_80; // @[AsyncQueue.scala 47:37]
  wire  _GEN_81; // @[AsyncQueue.scala 47:37]
  wire  _GEN_82; // @[AsyncQueue.scala 47:37]
  wire  _GEN_83; // @[AsyncQueue.scala 47:37]
  wire  _GEN_84; // @[AsyncQueue.scala 47:37]
  wire  _GEN_85; // @[AsyncQueue.scala 47:37]
  wire  _GEN_86; // @[AsyncQueue.scala 47:37]
  wire  _GEN_87; // @[AsyncQueue.scala 47:37]
  wire  _GEN_88; // @[AsyncQueue.scala 47:37]
  wire  _GEN_89; // @[AsyncQueue.scala 47:37]
  wire  _GEN_90; // @[AsyncQueue.scala 47:37]
  wire  _GEN_91; // @[AsyncQueue.scala 47:37]
  wire  _GEN_92; // @[AsyncQueue.scala 47:37]
  wire  _GEN_93; // @[AsyncQueue.scala 47:37]
  wire  _GEN_94; // @[AsyncQueue.scala 47:37]
  wire  _GEN_95; // @[AsyncQueue.scala 47:37]
  wire  _GEN_96; // @[AsyncQueue.scala 47:37]
  wire  _GEN_97; // @[AsyncQueue.scala 47:37]
  wire  _GEN_98; // @[AsyncQueue.scala 47:37]
  wire  _GEN_99; // @[AsyncQueue.scala 47:37]
  wire  _GEN_100; // @[AsyncQueue.scala 47:37]
  wire  _GEN_101; // @[AsyncQueue.scala 47:37]
  wire  _GEN_102; // @[AsyncQueue.scala 47:37]
  wire  _GEN_103; // @[AsyncQueue.scala 47:37]
  wire  _GEN_104; // @[AsyncQueue.scala 47:37]
  wire  _GEN_105; // @[AsyncQueue.scala 47:37]
  wire  _GEN_106; // @[AsyncQueue.scala 47:37]
  wire  _GEN_107; // @[AsyncQueue.scala 47:37]
  wire  _GEN_108; // @[AsyncQueue.scala 47:37]
  wire  _GEN_109; // @[AsyncQueue.scala 47:37]
  wire  _GEN_110; // @[AsyncQueue.scala 47:37]
  wire  _GEN_111; // @[AsyncQueue.scala 47:37]
  wire  _GEN_112; // @[AsyncQueue.scala 47:37]
  wire  _GEN_113; // @[AsyncQueue.scala 47:37]
  wire  _GEN_114; // @[AsyncQueue.scala 47:37]
  wire  _GEN_115; // @[AsyncQueue.scala 47:37]
  wire  _GEN_116; // @[AsyncQueue.scala 47:37]
  wire  _GEN_117; // @[AsyncQueue.scala 47:37]
  wire  _GEN_118; // @[AsyncQueue.scala 47:37]
  wire  _GEN_119; // @[AsyncQueue.scala 47:37]
  wire  _GEN_120; // @[AsyncQueue.scala 47:37]
  wire  _GEN_121; // @[AsyncQueue.scala 47:37]
  wire  _GEN_122; // @[AsyncQueue.scala 47:37]
  wire  _GEN_123; // @[AsyncQueue.scala 47:37]
  wire  _GEN_124; // @[AsyncQueue.scala 47:37]
  wire  _GEN_125; // @[AsyncQueue.scala 47:37]
  wire  _GEN_126; // @[AsyncQueue.scala 47:37]
  wire  _GEN_127; // @[AsyncQueue.scala 47:37]
  wire  _GEN_128; // @[AsyncQueue.scala 47:37]
  wire  _GEN_129; // @[AsyncQueue.scala 47:37]
  wire  _GEN_130; // @[AsyncQueue.scala 47:37]
  wire  _GEN_131; // @[AsyncQueue.scala 47:37]
  wire  _GEN_132; // @[AsyncQueue.scala 47:37]
  wire  _GEN_133; // @[AsyncQueue.scala 47:37]
  wire  _GEN_134; // @[AsyncQueue.scala 47:37]
  wire  _GEN_135; // @[AsyncQueue.scala 47:37]
  wire  _GEN_136; // @[AsyncQueue.scala 47:37]
  wire  _GEN_137; // @[AsyncQueue.scala 47:37]
  wire  _GEN_138; // @[AsyncQueue.scala 47:37]
  wire  _GEN_139; // @[AsyncQueue.scala 47:37]
  wire  _GEN_140; // @[AsyncQueue.scala 47:37]
  wire  _GEN_141; // @[AsyncQueue.scala 47:37]
  wire  _GEN_142; // @[AsyncQueue.scala 47:37]
  wire  _GEN_143; // @[AsyncQueue.scala 47:37]
  wire  _GEN_144; // @[AsyncQueue.scala 47:37]
  wire  _GEN_145; // @[AsyncQueue.scala 47:37]
  wire  _GEN_146; // @[AsyncQueue.scala 47:37]
  wire  _GEN_147; // @[AsyncQueue.scala 47:37]
  wire  _GEN_148; // @[AsyncQueue.scala 47:37]
  wire  _GEN_149; // @[AsyncQueue.scala 47:37]
  wire  _GEN_150; // @[AsyncQueue.scala 47:37]
  wire  _GEN_151; // @[AsyncQueue.scala 47:37]
  wire  _GEN_152; // @[AsyncQueue.scala 47:37]
  wire  _GEN_153; // @[AsyncQueue.scala 47:37]
  wire  _GEN_154; // @[AsyncQueue.scala 47:37]
  wire  _GEN_155; // @[AsyncQueue.scala 47:37]
  wire  _GEN_156; // @[AsyncQueue.scala 47:37]
  wire  _GEN_157; // @[AsyncQueue.scala 47:37]
  wire  _GEN_158; // @[AsyncQueue.scala 47:37]
  wire  _GEN_159; // @[AsyncQueue.scala 47:37]
  wire  _GEN_160; // @[AsyncQueue.scala 47:37]
  wire  _GEN_161; // @[AsyncQueue.scala 47:37]
  wire  _GEN_162; // @[AsyncQueue.scala 47:37]
  wire  _GEN_163; // @[AsyncQueue.scala 47:37]
  wire  _GEN_164; // @[AsyncQueue.scala 47:37]
  wire  _GEN_165; // @[AsyncQueue.scala 47:37]
  wire  _GEN_166; // @[AsyncQueue.scala 47:37]
  wire  _GEN_167; // @[AsyncQueue.scala 47:37]
  wire  _GEN_168; // @[AsyncQueue.scala 47:37]
  wire  _GEN_169; // @[AsyncQueue.scala 47:37]
  wire  _GEN_170; // @[AsyncQueue.scala 47:37]
  wire  _GEN_171; // @[AsyncQueue.scala 47:37]
  wire  _GEN_172; // @[AsyncQueue.scala 47:37]
  wire  _GEN_173; // @[AsyncQueue.scala 47:37]
  wire  _GEN_174; // @[AsyncQueue.scala 47:37]
  wire  _GEN_175; // @[AsyncQueue.scala 47:37]
  wire  _GEN_176; // @[AsyncQueue.scala 47:37]
  wire  _GEN_177; // @[AsyncQueue.scala 47:37]
  wire  _GEN_178; // @[AsyncQueue.scala 47:37]
  wire  _GEN_179; // @[AsyncQueue.scala 47:37]
  wire  _GEN_180; // @[AsyncQueue.scala 47:37]
  wire  _GEN_181; // @[AsyncQueue.scala 47:37]
  wire  _GEN_182; // @[AsyncQueue.scala 47:37]
  wire  _GEN_183; // @[AsyncQueue.scala 47:37]
  wire  _GEN_184; // @[AsyncQueue.scala 47:37]
  wire  _GEN_185; // @[AsyncQueue.scala 47:37]
  wire  _GEN_186; // @[AsyncQueue.scala 47:37]
  wire  _GEN_187; // @[AsyncQueue.scala 47:37]
  wire  _GEN_188; // @[AsyncQueue.scala 47:37]
  wire  _GEN_189; // @[AsyncQueue.scala 47:37]
  wire  _GEN_190; // @[AsyncQueue.scala 47:37]
  wire  _GEN_191; // @[AsyncQueue.scala 47:37]
  wire  _GEN_192; // @[AsyncQueue.scala 47:37]
  wire  _GEN_193; // @[AsyncQueue.scala 47:37]
  wire  _GEN_194; // @[AsyncQueue.scala 47:37]
  wire  _GEN_195; // @[AsyncQueue.scala 47:37]
  wire  _GEN_196; // @[AsyncQueue.scala 47:37]
  wire  _GEN_197; // @[AsyncQueue.scala 47:37]
  wire  _GEN_198; // @[AsyncQueue.scala 47:37]
  wire  _GEN_199; // @[AsyncQueue.scala 47:37]
  wire  _GEN_200; // @[AsyncQueue.scala 47:37]
  wire  _GEN_201; // @[AsyncQueue.scala 47:37]
  wire  _GEN_202; // @[AsyncQueue.scala 47:37]
  wire  _GEN_203; // @[AsyncQueue.scala 47:37]
  wire  _GEN_204; // @[AsyncQueue.scala 47:37]
  wire  _GEN_205; // @[AsyncQueue.scala 47:37]
  wire  _GEN_206; // @[AsyncQueue.scala 47:37]
  wire  _GEN_207; // @[AsyncQueue.scala 47:37]
  wire  _GEN_208; // @[AsyncQueue.scala 47:37]
  wire  _GEN_209; // @[AsyncQueue.scala 47:37]
  wire  _GEN_210; // @[AsyncQueue.scala 47:37]
  wire  _GEN_211; // @[AsyncQueue.scala 47:37]
  wire  _GEN_212; // @[AsyncQueue.scala 47:37]
  wire  _GEN_213; // @[AsyncQueue.scala 47:37]
  wire  _GEN_214; // @[AsyncQueue.scala 47:37]
  wire  _GEN_215; // @[AsyncQueue.scala 47:37]
  wire  _GEN_216; // @[AsyncQueue.scala 47:37]
  wire  _GEN_217; // @[AsyncQueue.scala 47:37]
  wire  _GEN_218; // @[AsyncQueue.scala 47:37]
  wire  _GEN_219; // @[AsyncQueue.scala 47:37]
  wire  _GEN_220; // @[AsyncQueue.scala 47:37]
  wire  _GEN_221; // @[AsyncQueue.scala 47:37]
  wire  _GEN_222; // @[AsyncQueue.scala 47:37]
  wire  _GEN_223; // @[AsyncQueue.scala 47:37]
  wire  _GEN_224; // @[AsyncQueue.scala 47:37]
  wire  _GEN_225; // @[AsyncQueue.scala 47:37]
  wire  _GEN_226; // @[AsyncQueue.scala 47:37]
  wire  _GEN_227; // @[AsyncQueue.scala 47:37]
  wire  _GEN_228; // @[AsyncQueue.scala 47:37]
  wire  _GEN_229; // @[AsyncQueue.scala 47:37]
  wire  _GEN_230; // @[AsyncQueue.scala 47:37]
  wire  _GEN_231; // @[AsyncQueue.scala 47:37]
  wire  _GEN_232; // @[AsyncQueue.scala 47:37]
  wire  _GEN_233; // @[AsyncQueue.scala 47:37]
  wire  _GEN_234; // @[AsyncQueue.scala 47:37]
  wire  _GEN_235; // @[AsyncQueue.scala 47:37]
  wire  _GEN_236; // @[AsyncQueue.scala 47:37]
  wire  _GEN_237; // @[AsyncQueue.scala 47:37]
  wire  _GEN_238; // @[AsyncQueue.scala 47:37]
  wire  _GEN_239; // @[AsyncQueue.scala 47:37]
  wire  _GEN_240; // @[AsyncQueue.scala 47:37]
  wire  _GEN_241; // @[AsyncQueue.scala 47:37]
  wire  _GEN_242; // @[AsyncQueue.scala 47:37]
  wire  _GEN_243; // @[AsyncQueue.scala 47:37]
  wire  _GEN_244; // @[AsyncQueue.scala 47:37]
  wire  _GEN_245; // @[AsyncQueue.scala 47:37]
  wire  _GEN_246; // @[AsyncQueue.scala 47:37]
  wire  _GEN_247; // @[AsyncQueue.scala 47:37]
  wire  _GEN_248; // @[AsyncQueue.scala 47:37]
  wire  _GEN_249; // @[AsyncQueue.scala 47:37]
  wire  _GEN_250; // @[AsyncQueue.scala 47:37]
  wire  _GEN_251; // @[AsyncQueue.scala 47:37]
  wire  _GEN_252; // @[AsyncQueue.scala 47:37]
  wire  _GEN_253; // @[AsyncQueue.scala 47:37]
  wire  _GEN_254; // @[AsyncQueue.scala 47:37]
  wire  _GEN_255; // @[AsyncQueue.scala 47:37]
  wire  _GEN_256; // @[AsyncQueue.scala 47:37]
  wire  _GEN_257; // @[AsyncQueue.scala 47:24]
  wire  _GEN_258; // @[AsyncQueue.scala 47:24]
  wire  _GEN_259; // @[AsyncQueue.scala 47:24]
  wire  _GEN_260; // @[AsyncQueue.scala 47:24]
  wire  _GEN_261; // @[AsyncQueue.scala 47:24]
  wire  _GEN_262; // @[AsyncQueue.scala 47:24]
  wire  _GEN_263; // @[AsyncQueue.scala 47:24]
  wire  _GEN_264; // @[AsyncQueue.scala 47:24]
  wire  _GEN_265; // @[AsyncQueue.scala 47:24]
  wire  _GEN_266; // @[AsyncQueue.scala 47:24]
  wire  _GEN_267; // @[AsyncQueue.scala 47:24]
  wire  _GEN_268; // @[AsyncQueue.scala 47:24]
  wire  _GEN_269; // @[AsyncQueue.scala 47:24]
  wire  _GEN_270; // @[AsyncQueue.scala 47:24]
  wire  _GEN_271; // @[AsyncQueue.scala 47:24]
  wire  _GEN_272; // @[AsyncQueue.scala 47:24]
  wire  _GEN_273; // @[AsyncQueue.scala 47:24]
  wire  _GEN_274; // @[AsyncQueue.scala 47:24]
  wire  _GEN_275; // @[AsyncQueue.scala 47:24]
  wire  _GEN_276; // @[AsyncQueue.scala 47:24]
  wire  _GEN_277; // @[AsyncQueue.scala 47:24]
  wire  _GEN_278; // @[AsyncQueue.scala 47:24]
  wire  _GEN_279; // @[AsyncQueue.scala 47:24]
  wire  _GEN_280; // @[AsyncQueue.scala 47:24]
  wire  _GEN_281; // @[AsyncQueue.scala 47:24]
  wire  _GEN_282; // @[AsyncQueue.scala 47:24]
  wire  _GEN_283; // @[AsyncQueue.scala 47:24]
  wire  _GEN_284; // @[AsyncQueue.scala 47:24]
  wire  _GEN_285; // @[AsyncQueue.scala 47:24]
  wire  _GEN_286; // @[AsyncQueue.scala 47:24]
  wire  _GEN_287; // @[AsyncQueue.scala 47:24]
  wire  _GEN_288; // @[AsyncQueue.scala 47:24]
  wire  _GEN_289; // @[AsyncQueue.scala 47:24]
  wire  _GEN_290; // @[AsyncQueue.scala 47:24]
  wire  _GEN_291; // @[AsyncQueue.scala 47:24]
  wire  _GEN_292; // @[AsyncQueue.scala 47:24]
  wire  _GEN_293; // @[AsyncQueue.scala 47:24]
  wire  _GEN_294; // @[AsyncQueue.scala 47:24]
  wire  _GEN_295; // @[AsyncQueue.scala 47:24]
  wire  _GEN_296; // @[AsyncQueue.scala 47:24]
  wire  _GEN_297; // @[AsyncQueue.scala 47:24]
  wire  _GEN_298; // @[AsyncQueue.scala 47:24]
  wire  _GEN_299; // @[AsyncQueue.scala 47:24]
  wire  _GEN_300; // @[AsyncQueue.scala 47:24]
  wire  _GEN_301; // @[AsyncQueue.scala 47:24]
  wire  _GEN_302; // @[AsyncQueue.scala 47:24]
  wire  _GEN_303; // @[AsyncQueue.scala 47:24]
  wire  _GEN_304; // @[AsyncQueue.scala 47:24]
  wire  _GEN_305; // @[AsyncQueue.scala 47:24]
  wire  _GEN_306; // @[AsyncQueue.scala 47:24]
  wire  _GEN_307; // @[AsyncQueue.scala 47:24]
  wire  _GEN_308; // @[AsyncQueue.scala 47:24]
  wire  _GEN_309; // @[AsyncQueue.scala 47:24]
  wire  _GEN_310; // @[AsyncQueue.scala 47:24]
  wire  _GEN_311; // @[AsyncQueue.scala 47:24]
  wire  _GEN_312; // @[AsyncQueue.scala 47:24]
  wire  _GEN_313; // @[AsyncQueue.scala 47:24]
  wire  _GEN_314; // @[AsyncQueue.scala 47:24]
  wire  _GEN_315; // @[AsyncQueue.scala 47:24]
  wire  _GEN_316; // @[AsyncQueue.scala 47:24]
  wire  _GEN_317; // @[AsyncQueue.scala 47:24]
  wire  _GEN_318; // @[AsyncQueue.scala 47:24]
  wire  _GEN_319; // @[AsyncQueue.scala 47:24]
  wire  _GEN_320; // @[AsyncQueue.scala 47:24]
  wire  _GEN_321; // @[AsyncQueue.scala 47:24]
  wire  _GEN_322; // @[AsyncQueue.scala 47:24]
  wire  _GEN_323; // @[AsyncQueue.scala 47:24]
  wire  _GEN_324; // @[AsyncQueue.scala 47:24]
  wire  _GEN_325; // @[AsyncQueue.scala 47:24]
  wire  _GEN_326; // @[AsyncQueue.scala 47:24]
  wire  _GEN_327; // @[AsyncQueue.scala 47:24]
  wire  _GEN_328; // @[AsyncQueue.scala 47:24]
  wire  _GEN_329; // @[AsyncQueue.scala 47:24]
  wire  _GEN_330; // @[AsyncQueue.scala 47:24]
  wire  _GEN_331; // @[AsyncQueue.scala 47:24]
  wire  _GEN_332; // @[AsyncQueue.scala 47:24]
  wire  _GEN_333; // @[AsyncQueue.scala 47:24]
  wire  _GEN_334; // @[AsyncQueue.scala 47:24]
  wire  _GEN_335; // @[AsyncQueue.scala 47:24]
  wire  _GEN_336; // @[AsyncQueue.scala 47:24]
  wire  _GEN_337; // @[AsyncQueue.scala 47:24]
  wire  _GEN_338; // @[AsyncQueue.scala 47:24]
  wire  _GEN_339; // @[AsyncQueue.scala 47:24]
  wire  _GEN_340; // @[AsyncQueue.scala 47:24]
  wire  _GEN_341; // @[AsyncQueue.scala 47:24]
  wire  _GEN_342; // @[AsyncQueue.scala 47:24]
  wire  _GEN_343; // @[AsyncQueue.scala 47:24]
  wire  _GEN_344; // @[AsyncQueue.scala 47:24]
  wire  _GEN_345; // @[AsyncQueue.scala 47:24]
  wire  _GEN_346; // @[AsyncQueue.scala 47:24]
  wire  _GEN_347; // @[AsyncQueue.scala 47:24]
  wire  _GEN_348; // @[AsyncQueue.scala 47:24]
  wire  _GEN_349; // @[AsyncQueue.scala 47:24]
  wire  _GEN_350; // @[AsyncQueue.scala 47:24]
  wire  _GEN_351; // @[AsyncQueue.scala 47:24]
  wire  _GEN_352; // @[AsyncQueue.scala 47:24]
  wire  _GEN_353; // @[AsyncQueue.scala 47:24]
  wire  _GEN_354; // @[AsyncQueue.scala 47:24]
  wire  _GEN_355; // @[AsyncQueue.scala 47:24]
  wire  _GEN_356; // @[AsyncQueue.scala 47:24]
  wire  _GEN_357; // @[AsyncQueue.scala 47:24]
  wire  _GEN_358; // @[AsyncQueue.scala 47:24]
  wire  _GEN_359; // @[AsyncQueue.scala 47:24]
  wire  _GEN_360; // @[AsyncQueue.scala 47:24]
  wire  _GEN_361; // @[AsyncQueue.scala 47:24]
  wire  _GEN_362; // @[AsyncQueue.scala 47:24]
  wire  _GEN_363; // @[AsyncQueue.scala 47:24]
  wire  _GEN_364; // @[AsyncQueue.scala 47:24]
  wire  _GEN_365; // @[AsyncQueue.scala 47:24]
  wire  _GEN_366; // @[AsyncQueue.scala 47:24]
  wire  _GEN_367; // @[AsyncQueue.scala 47:24]
  wire  _GEN_368; // @[AsyncQueue.scala 47:24]
  wire  _GEN_369; // @[AsyncQueue.scala 47:24]
  wire  _GEN_370; // @[AsyncQueue.scala 47:24]
  wire  _GEN_371; // @[AsyncQueue.scala 47:24]
  wire  _GEN_372; // @[AsyncQueue.scala 47:24]
  wire  _GEN_373; // @[AsyncQueue.scala 47:24]
  wire  _GEN_374; // @[AsyncQueue.scala 47:24]
  wire  _GEN_375; // @[AsyncQueue.scala 47:24]
  wire  _GEN_376; // @[AsyncQueue.scala 47:24]
  wire  _GEN_377; // @[AsyncQueue.scala 47:24]
  wire  _GEN_378; // @[AsyncQueue.scala 47:24]
  wire  _GEN_379; // @[AsyncQueue.scala 47:24]
  wire  _GEN_380; // @[AsyncQueue.scala 47:24]
  wire  _GEN_381; // @[AsyncQueue.scala 47:24]
  wire  _GEN_382; // @[AsyncQueue.scala 47:24]
  wire  _GEN_383; // @[AsyncQueue.scala 47:24]
  wire  _GEN_384; // @[AsyncQueue.scala 47:24]
  wire  _GEN_385; // @[AsyncQueue.scala 47:24]
  wire  _GEN_386; // @[AsyncQueue.scala 47:24]
  wire  _GEN_387; // @[AsyncQueue.scala 47:24]
  wire  _GEN_388; // @[AsyncQueue.scala 47:24]
  wire  _GEN_389; // @[AsyncQueue.scala 47:24]
  wire  _GEN_390; // @[AsyncQueue.scala 47:24]
  wire  _GEN_391; // @[AsyncQueue.scala 47:24]
  wire  _GEN_392; // @[AsyncQueue.scala 47:24]
  wire  _GEN_393; // @[AsyncQueue.scala 47:24]
  wire  _GEN_394; // @[AsyncQueue.scala 47:24]
  wire  _GEN_395; // @[AsyncQueue.scala 47:24]
  wire  _GEN_396; // @[AsyncQueue.scala 47:24]
  wire  _GEN_397; // @[AsyncQueue.scala 47:24]
  wire  _GEN_398; // @[AsyncQueue.scala 47:24]
  wire  _GEN_399; // @[AsyncQueue.scala 47:24]
  wire  _GEN_400; // @[AsyncQueue.scala 47:24]
  wire  _GEN_401; // @[AsyncQueue.scala 47:24]
  wire  _GEN_402; // @[AsyncQueue.scala 47:24]
  wire  _GEN_403; // @[AsyncQueue.scala 47:24]
  wire  _GEN_404; // @[AsyncQueue.scala 47:24]
  wire  _GEN_405; // @[AsyncQueue.scala 47:24]
  wire  _GEN_406; // @[AsyncQueue.scala 47:24]
  wire  _GEN_407; // @[AsyncQueue.scala 47:24]
  wire  _GEN_408; // @[AsyncQueue.scala 47:24]
  wire  _GEN_409; // @[AsyncQueue.scala 47:24]
  wire  _GEN_410; // @[AsyncQueue.scala 47:24]
  wire  _GEN_411; // @[AsyncQueue.scala 47:24]
  wire  _GEN_412; // @[AsyncQueue.scala 47:24]
  wire  _GEN_413; // @[AsyncQueue.scala 47:24]
  wire  _GEN_414; // @[AsyncQueue.scala 47:24]
  wire  _GEN_415; // @[AsyncQueue.scala 47:24]
  wire  _GEN_416; // @[AsyncQueue.scala 47:24]
  wire  _GEN_417; // @[AsyncQueue.scala 47:24]
  wire  _GEN_418; // @[AsyncQueue.scala 47:24]
  wire  _GEN_419; // @[AsyncQueue.scala 47:24]
  wire  _GEN_420; // @[AsyncQueue.scala 47:24]
  wire  _GEN_421; // @[AsyncQueue.scala 47:24]
  wire  _GEN_422; // @[AsyncQueue.scala 47:24]
  wire  _GEN_423; // @[AsyncQueue.scala 47:24]
  wire  _GEN_424; // @[AsyncQueue.scala 47:24]
  wire  _GEN_425; // @[AsyncQueue.scala 47:24]
  wire  _GEN_426; // @[AsyncQueue.scala 47:24]
  wire  _GEN_427; // @[AsyncQueue.scala 47:24]
  wire  _GEN_428; // @[AsyncQueue.scala 47:24]
  wire  _GEN_429; // @[AsyncQueue.scala 47:24]
  wire  _GEN_430; // @[AsyncQueue.scala 47:24]
  wire  _GEN_431; // @[AsyncQueue.scala 47:24]
  wire  _GEN_432; // @[AsyncQueue.scala 47:24]
  wire  _GEN_433; // @[AsyncQueue.scala 47:24]
  wire  _GEN_434; // @[AsyncQueue.scala 47:24]
  wire  _GEN_435; // @[AsyncQueue.scala 47:24]
  wire  _GEN_436; // @[AsyncQueue.scala 47:24]
  wire  _GEN_437; // @[AsyncQueue.scala 47:24]
  wire  _GEN_438; // @[AsyncQueue.scala 47:24]
  wire  _GEN_439; // @[AsyncQueue.scala 47:24]
  wire  _GEN_440; // @[AsyncQueue.scala 47:24]
  wire  _GEN_441; // @[AsyncQueue.scala 47:24]
  wire  _GEN_442; // @[AsyncQueue.scala 47:24]
  wire  _GEN_443; // @[AsyncQueue.scala 47:24]
  wire  _GEN_444; // @[AsyncQueue.scala 47:24]
  wire  _GEN_445; // @[AsyncQueue.scala 47:24]
  wire  _GEN_446; // @[AsyncQueue.scala 47:24]
  wire  _GEN_447; // @[AsyncQueue.scala 47:24]
  wire  _GEN_448; // @[AsyncQueue.scala 47:24]
  wire  _GEN_449; // @[AsyncQueue.scala 47:24]
  wire  _GEN_450; // @[AsyncQueue.scala 47:24]
  wire  _GEN_451; // @[AsyncQueue.scala 47:24]
  wire  _GEN_452; // @[AsyncQueue.scala 47:24]
  wire  _GEN_453; // @[AsyncQueue.scala 47:24]
  wire  _GEN_454; // @[AsyncQueue.scala 47:24]
  wire  _GEN_455; // @[AsyncQueue.scala 47:24]
  wire  _GEN_456; // @[AsyncQueue.scala 47:24]
  wire  _GEN_457; // @[AsyncQueue.scala 47:24]
  wire  _GEN_458; // @[AsyncQueue.scala 47:24]
  wire  _GEN_459; // @[AsyncQueue.scala 47:24]
  wire  _GEN_460; // @[AsyncQueue.scala 47:24]
  wire  _GEN_461; // @[AsyncQueue.scala 47:24]
  wire  _GEN_462; // @[AsyncQueue.scala 47:24]
  wire  _GEN_463; // @[AsyncQueue.scala 47:24]
  wire  _GEN_464; // @[AsyncQueue.scala 47:24]
  wire  _GEN_465; // @[AsyncQueue.scala 47:24]
  wire  _GEN_466; // @[AsyncQueue.scala 47:24]
  wire  _GEN_467; // @[AsyncQueue.scala 47:24]
  wire  _GEN_468; // @[AsyncQueue.scala 47:24]
  wire  _GEN_469; // @[AsyncQueue.scala 47:24]
  wire  _GEN_470; // @[AsyncQueue.scala 47:24]
  wire  _GEN_471; // @[AsyncQueue.scala 47:24]
  wire  _GEN_472; // @[AsyncQueue.scala 47:24]
  wire  _GEN_473; // @[AsyncQueue.scala 47:24]
  wire  _GEN_474; // @[AsyncQueue.scala 47:24]
  wire  _GEN_475; // @[AsyncQueue.scala 47:24]
  wire  _GEN_476; // @[AsyncQueue.scala 47:24]
  wire  _GEN_477; // @[AsyncQueue.scala 47:24]
  wire  _GEN_478; // @[AsyncQueue.scala 47:24]
  wire  _GEN_479; // @[AsyncQueue.scala 47:24]
  wire  _GEN_480; // @[AsyncQueue.scala 47:24]
  wire  _GEN_481; // @[AsyncQueue.scala 47:24]
  wire  _GEN_482; // @[AsyncQueue.scala 47:24]
  wire  _GEN_483; // @[AsyncQueue.scala 47:24]
  wire  _GEN_484; // @[AsyncQueue.scala 47:24]
  wire  _GEN_485; // @[AsyncQueue.scala 47:24]
  wire  _GEN_486; // @[AsyncQueue.scala 47:24]
  wire  _GEN_487; // @[AsyncQueue.scala 47:24]
  wire  _GEN_488; // @[AsyncQueue.scala 47:24]
  wire  _GEN_489; // @[AsyncQueue.scala 47:24]
  wire  _GEN_490; // @[AsyncQueue.scala 47:24]
  wire  _GEN_491; // @[AsyncQueue.scala 47:24]
  wire  _GEN_492; // @[AsyncQueue.scala 47:24]
  wire  _GEN_493; // @[AsyncQueue.scala 47:24]
  wire  _GEN_494; // @[AsyncQueue.scala 47:24]
  wire  _GEN_495; // @[AsyncQueue.scala 47:24]
  wire  _GEN_496; // @[AsyncQueue.scala 47:24]
  wire  _GEN_497; // @[AsyncQueue.scala 47:24]
  wire  _GEN_498; // @[AsyncQueue.scala 47:24]
  wire  _GEN_499; // @[AsyncQueue.scala 47:24]
  wire  _GEN_500; // @[AsyncQueue.scala 47:24]
  wire  _GEN_501; // @[AsyncQueue.scala 47:24]
  wire  _GEN_502; // @[AsyncQueue.scala 47:24]
  wire  _GEN_503; // @[AsyncQueue.scala 47:24]
  wire  _GEN_504; // @[AsyncQueue.scala 47:24]
  wire  _GEN_505; // @[AsyncQueue.scala 47:24]
  wire  _GEN_506; // @[AsyncQueue.scala 47:24]
  wire  _GEN_507; // @[AsyncQueue.scala 47:24]
  wire  _GEN_508; // @[AsyncQueue.scala 47:24]
  wire  _GEN_509; // @[AsyncQueue.scala 47:24]
  wire  _GEN_510; // @[AsyncQueue.scala 47:24]
  wire  _GEN_511; // @[AsyncQueue.scala 47:24]
  wire  _GEN_512; // @[AsyncQueue.scala 47:24]
  wire  ready_reg_1; // @[AsyncQueue.scala 49:59]
  wire  _T_558; // @[AsyncQueue.scala 50:29]
  wire  _T_563; // @[AsyncQueue.scala 62:36]
  wire  _T_564; // @[AsyncQueue.scala 62:33]
  AsyncResetRegVec_w9_i0 widx_bin ( // @[AsyncResetReg.scala 110:21]
    .clock(widx_bin_clock),
    .reset(widx_bin_reset),
    .io_d(widx_bin_io_d),
    .io_q(widx_bin_io_q),
    .io_en(widx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w9_d3_i0 ridx_gray ( // @[ShiftReg.scala 47:23]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q)
  );
  AsyncResetRegVec_w1_i0 ready_reg ( // @[AsyncResetReg.scala 110:21]
    .clock(ready_reg_clock),
    .reset(ready_reg_reset),
    .io_d(ready_reg_io_d),
    .io_q(ready_reg_io_q),
    .io_en(ready_reg_io_en)
  );
  AsyncResetRegVec_w9_i0 widx_gray ( // @[AsyncResetReg.scala 110:21]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q),
    .io_en(widx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 59:30]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 ( // @[AsyncQueue.scala 60:30]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 ( // @[AsyncQueue.scala 61:30]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  assign _T_536 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 30:37]
  assign sink_ready = AsyncValidSync_2_io_out;
  assign _T_538 = sink_ready == 1'h0; // @[AsyncQueue.scala 42:49]
  assign _GEN_513 = {{8'd0}, _T_536}; // @[AsyncQueue.scala 11:47]
  assign _T_543 = widx_bin_io_q + _GEN_513; // @[AsyncQueue.scala 11:47]
  assign _T_544 = _T_543[8:0]; // @[AsyncQueue.scala 11:47]
  assign _T_545 = _T_538 ? 9'h0 : _T_544; // @[AsyncQueue.scala 11:23]
  assign _T_547 = _T_545 >> 1'h1; // @[AsyncQueue.scala 12:32]
  assign widx = _T_545 ^ _T_547; // @[AsyncQueue.scala 12:17]
  assign ridx = ridx_gray_io_q; // @[ShiftReg.scala 50:24]
  assign _T_550 = ridx ^ 9'h180; // @[AsyncQueue.scala 44:44]
  assign _T_551 = widx != _T_550; // @[AsyncQueue.scala 44:34]
  assign ready = sink_ready & _T_551; // @[AsyncQueue.scala 44:26]
  assign _T_552 = io_widx[7:0]; // @[AsyncQueue.scala 46:51]
  assign _T_553 = io_widx[8]; // @[AsyncQueue.scala 46:73]
  assign _GEN_514 = {{7'd0}, _T_553}; // @[AsyncQueue.scala 46:86]
  assign _T_554 = _GEN_514 << 7; // @[AsyncQueue.scala 46:86]
  assign index = _T_552 ^ _T_554; // @[AsyncQueue.scala 46:63]
  assign _GEN_1 = 8'h0 == index ? io_enq_bits : mem_0; // @[AsyncQueue.scala 47:37]
  assign _GEN_2 = 8'h1 == index ? io_enq_bits : mem_1; // @[AsyncQueue.scala 47:37]
  assign _GEN_3 = 8'h2 == index ? io_enq_bits : mem_2; // @[AsyncQueue.scala 47:37]
  assign _GEN_4 = 8'h3 == index ? io_enq_bits : mem_3; // @[AsyncQueue.scala 47:37]
  assign _GEN_5 = 8'h4 == index ? io_enq_bits : mem_4; // @[AsyncQueue.scala 47:37]
  assign _GEN_6 = 8'h5 == index ? io_enq_bits : mem_5; // @[AsyncQueue.scala 47:37]
  assign _GEN_7 = 8'h6 == index ? io_enq_bits : mem_6; // @[AsyncQueue.scala 47:37]
  assign _GEN_8 = 8'h7 == index ? io_enq_bits : mem_7; // @[AsyncQueue.scala 47:37]
  assign _GEN_9 = 8'h8 == index ? io_enq_bits : mem_8; // @[AsyncQueue.scala 47:37]
  assign _GEN_10 = 8'h9 == index ? io_enq_bits : mem_9; // @[AsyncQueue.scala 47:37]
  assign _GEN_11 = 8'ha == index ? io_enq_bits : mem_10; // @[AsyncQueue.scala 47:37]
  assign _GEN_12 = 8'hb == index ? io_enq_bits : mem_11; // @[AsyncQueue.scala 47:37]
  assign _GEN_13 = 8'hc == index ? io_enq_bits : mem_12; // @[AsyncQueue.scala 47:37]
  assign _GEN_14 = 8'hd == index ? io_enq_bits : mem_13; // @[AsyncQueue.scala 47:37]
  assign _GEN_15 = 8'he == index ? io_enq_bits : mem_14; // @[AsyncQueue.scala 47:37]
  assign _GEN_16 = 8'hf == index ? io_enq_bits : mem_15; // @[AsyncQueue.scala 47:37]
  assign _GEN_17 = 8'h10 == index ? io_enq_bits : mem_16; // @[AsyncQueue.scala 47:37]
  assign _GEN_18 = 8'h11 == index ? io_enq_bits : mem_17; // @[AsyncQueue.scala 47:37]
  assign _GEN_19 = 8'h12 == index ? io_enq_bits : mem_18; // @[AsyncQueue.scala 47:37]
  assign _GEN_20 = 8'h13 == index ? io_enq_bits : mem_19; // @[AsyncQueue.scala 47:37]
  assign _GEN_21 = 8'h14 == index ? io_enq_bits : mem_20; // @[AsyncQueue.scala 47:37]
  assign _GEN_22 = 8'h15 == index ? io_enq_bits : mem_21; // @[AsyncQueue.scala 47:37]
  assign _GEN_23 = 8'h16 == index ? io_enq_bits : mem_22; // @[AsyncQueue.scala 47:37]
  assign _GEN_24 = 8'h17 == index ? io_enq_bits : mem_23; // @[AsyncQueue.scala 47:37]
  assign _GEN_25 = 8'h18 == index ? io_enq_bits : mem_24; // @[AsyncQueue.scala 47:37]
  assign _GEN_26 = 8'h19 == index ? io_enq_bits : mem_25; // @[AsyncQueue.scala 47:37]
  assign _GEN_27 = 8'h1a == index ? io_enq_bits : mem_26; // @[AsyncQueue.scala 47:37]
  assign _GEN_28 = 8'h1b == index ? io_enq_bits : mem_27; // @[AsyncQueue.scala 47:37]
  assign _GEN_29 = 8'h1c == index ? io_enq_bits : mem_28; // @[AsyncQueue.scala 47:37]
  assign _GEN_30 = 8'h1d == index ? io_enq_bits : mem_29; // @[AsyncQueue.scala 47:37]
  assign _GEN_31 = 8'h1e == index ? io_enq_bits : mem_30; // @[AsyncQueue.scala 47:37]
  assign _GEN_32 = 8'h1f == index ? io_enq_bits : mem_31; // @[AsyncQueue.scala 47:37]
  assign _GEN_33 = 8'h20 == index ? io_enq_bits : mem_32; // @[AsyncQueue.scala 47:37]
  assign _GEN_34 = 8'h21 == index ? io_enq_bits : mem_33; // @[AsyncQueue.scala 47:37]
  assign _GEN_35 = 8'h22 == index ? io_enq_bits : mem_34; // @[AsyncQueue.scala 47:37]
  assign _GEN_36 = 8'h23 == index ? io_enq_bits : mem_35; // @[AsyncQueue.scala 47:37]
  assign _GEN_37 = 8'h24 == index ? io_enq_bits : mem_36; // @[AsyncQueue.scala 47:37]
  assign _GEN_38 = 8'h25 == index ? io_enq_bits : mem_37; // @[AsyncQueue.scala 47:37]
  assign _GEN_39 = 8'h26 == index ? io_enq_bits : mem_38; // @[AsyncQueue.scala 47:37]
  assign _GEN_40 = 8'h27 == index ? io_enq_bits : mem_39; // @[AsyncQueue.scala 47:37]
  assign _GEN_41 = 8'h28 == index ? io_enq_bits : mem_40; // @[AsyncQueue.scala 47:37]
  assign _GEN_42 = 8'h29 == index ? io_enq_bits : mem_41; // @[AsyncQueue.scala 47:37]
  assign _GEN_43 = 8'h2a == index ? io_enq_bits : mem_42; // @[AsyncQueue.scala 47:37]
  assign _GEN_44 = 8'h2b == index ? io_enq_bits : mem_43; // @[AsyncQueue.scala 47:37]
  assign _GEN_45 = 8'h2c == index ? io_enq_bits : mem_44; // @[AsyncQueue.scala 47:37]
  assign _GEN_46 = 8'h2d == index ? io_enq_bits : mem_45; // @[AsyncQueue.scala 47:37]
  assign _GEN_47 = 8'h2e == index ? io_enq_bits : mem_46; // @[AsyncQueue.scala 47:37]
  assign _GEN_48 = 8'h2f == index ? io_enq_bits : mem_47; // @[AsyncQueue.scala 47:37]
  assign _GEN_49 = 8'h30 == index ? io_enq_bits : mem_48; // @[AsyncQueue.scala 47:37]
  assign _GEN_50 = 8'h31 == index ? io_enq_bits : mem_49; // @[AsyncQueue.scala 47:37]
  assign _GEN_51 = 8'h32 == index ? io_enq_bits : mem_50; // @[AsyncQueue.scala 47:37]
  assign _GEN_52 = 8'h33 == index ? io_enq_bits : mem_51; // @[AsyncQueue.scala 47:37]
  assign _GEN_53 = 8'h34 == index ? io_enq_bits : mem_52; // @[AsyncQueue.scala 47:37]
  assign _GEN_54 = 8'h35 == index ? io_enq_bits : mem_53; // @[AsyncQueue.scala 47:37]
  assign _GEN_55 = 8'h36 == index ? io_enq_bits : mem_54; // @[AsyncQueue.scala 47:37]
  assign _GEN_56 = 8'h37 == index ? io_enq_bits : mem_55; // @[AsyncQueue.scala 47:37]
  assign _GEN_57 = 8'h38 == index ? io_enq_bits : mem_56; // @[AsyncQueue.scala 47:37]
  assign _GEN_58 = 8'h39 == index ? io_enq_bits : mem_57; // @[AsyncQueue.scala 47:37]
  assign _GEN_59 = 8'h3a == index ? io_enq_bits : mem_58; // @[AsyncQueue.scala 47:37]
  assign _GEN_60 = 8'h3b == index ? io_enq_bits : mem_59; // @[AsyncQueue.scala 47:37]
  assign _GEN_61 = 8'h3c == index ? io_enq_bits : mem_60; // @[AsyncQueue.scala 47:37]
  assign _GEN_62 = 8'h3d == index ? io_enq_bits : mem_61; // @[AsyncQueue.scala 47:37]
  assign _GEN_63 = 8'h3e == index ? io_enq_bits : mem_62; // @[AsyncQueue.scala 47:37]
  assign _GEN_64 = 8'h3f == index ? io_enq_bits : mem_63; // @[AsyncQueue.scala 47:37]
  assign _GEN_65 = 8'h40 == index ? io_enq_bits : mem_64; // @[AsyncQueue.scala 47:37]
  assign _GEN_66 = 8'h41 == index ? io_enq_bits : mem_65; // @[AsyncQueue.scala 47:37]
  assign _GEN_67 = 8'h42 == index ? io_enq_bits : mem_66; // @[AsyncQueue.scala 47:37]
  assign _GEN_68 = 8'h43 == index ? io_enq_bits : mem_67; // @[AsyncQueue.scala 47:37]
  assign _GEN_69 = 8'h44 == index ? io_enq_bits : mem_68; // @[AsyncQueue.scala 47:37]
  assign _GEN_70 = 8'h45 == index ? io_enq_bits : mem_69; // @[AsyncQueue.scala 47:37]
  assign _GEN_71 = 8'h46 == index ? io_enq_bits : mem_70; // @[AsyncQueue.scala 47:37]
  assign _GEN_72 = 8'h47 == index ? io_enq_bits : mem_71; // @[AsyncQueue.scala 47:37]
  assign _GEN_73 = 8'h48 == index ? io_enq_bits : mem_72; // @[AsyncQueue.scala 47:37]
  assign _GEN_74 = 8'h49 == index ? io_enq_bits : mem_73; // @[AsyncQueue.scala 47:37]
  assign _GEN_75 = 8'h4a == index ? io_enq_bits : mem_74; // @[AsyncQueue.scala 47:37]
  assign _GEN_76 = 8'h4b == index ? io_enq_bits : mem_75; // @[AsyncQueue.scala 47:37]
  assign _GEN_77 = 8'h4c == index ? io_enq_bits : mem_76; // @[AsyncQueue.scala 47:37]
  assign _GEN_78 = 8'h4d == index ? io_enq_bits : mem_77; // @[AsyncQueue.scala 47:37]
  assign _GEN_79 = 8'h4e == index ? io_enq_bits : mem_78; // @[AsyncQueue.scala 47:37]
  assign _GEN_80 = 8'h4f == index ? io_enq_bits : mem_79; // @[AsyncQueue.scala 47:37]
  assign _GEN_81 = 8'h50 == index ? io_enq_bits : mem_80; // @[AsyncQueue.scala 47:37]
  assign _GEN_82 = 8'h51 == index ? io_enq_bits : mem_81; // @[AsyncQueue.scala 47:37]
  assign _GEN_83 = 8'h52 == index ? io_enq_bits : mem_82; // @[AsyncQueue.scala 47:37]
  assign _GEN_84 = 8'h53 == index ? io_enq_bits : mem_83; // @[AsyncQueue.scala 47:37]
  assign _GEN_85 = 8'h54 == index ? io_enq_bits : mem_84; // @[AsyncQueue.scala 47:37]
  assign _GEN_86 = 8'h55 == index ? io_enq_bits : mem_85; // @[AsyncQueue.scala 47:37]
  assign _GEN_87 = 8'h56 == index ? io_enq_bits : mem_86; // @[AsyncQueue.scala 47:37]
  assign _GEN_88 = 8'h57 == index ? io_enq_bits : mem_87; // @[AsyncQueue.scala 47:37]
  assign _GEN_89 = 8'h58 == index ? io_enq_bits : mem_88; // @[AsyncQueue.scala 47:37]
  assign _GEN_90 = 8'h59 == index ? io_enq_bits : mem_89; // @[AsyncQueue.scala 47:37]
  assign _GEN_91 = 8'h5a == index ? io_enq_bits : mem_90; // @[AsyncQueue.scala 47:37]
  assign _GEN_92 = 8'h5b == index ? io_enq_bits : mem_91; // @[AsyncQueue.scala 47:37]
  assign _GEN_93 = 8'h5c == index ? io_enq_bits : mem_92; // @[AsyncQueue.scala 47:37]
  assign _GEN_94 = 8'h5d == index ? io_enq_bits : mem_93; // @[AsyncQueue.scala 47:37]
  assign _GEN_95 = 8'h5e == index ? io_enq_bits : mem_94; // @[AsyncQueue.scala 47:37]
  assign _GEN_96 = 8'h5f == index ? io_enq_bits : mem_95; // @[AsyncQueue.scala 47:37]
  assign _GEN_97 = 8'h60 == index ? io_enq_bits : mem_96; // @[AsyncQueue.scala 47:37]
  assign _GEN_98 = 8'h61 == index ? io_enq_bits : mem_97; // @[AsyncQueue.scala 47:37]
  assign _GEN_99 = 8'h62 == index ? io_enq_bits : mem_98; // @[AsyncQueue.scala 47:37]
  assign _GEN_100 = 8'h63 == index ? io_enq_bits : mem_99; // @[AsyncQueue.scala 47:37]
  assign _GEN_101 = 8'h64 == index ? io_enq_bits : mem_100; // @[AsyncQueue.scala 47:37]
  assign _GEN_102 = 8'h65 == index ? io_enq_bits : mem_101; // @[AsyncQueue.scala 47:37]
  assign _GEN_103 = 8'h66 == index ? io_enq_bits : mem_102; // @[AsyncQueue.scala 47:37]
  assign _GEN_104 = 8'h67 == index ? io_enq_bits : mem_103; // @[AsyncQueue.scala 47:37]
  assign _GEN_105 = 8'h68 == index ? io_enq_bits : mem_104; // @[AsyncQueue.scala 47:37]
  assign _GEN_106 = 8'h69 == index ? io_enq_bits : mem_105; // @[AsyncQueue.scala 47:37]
  assign _GEN_107 = 8'h6a == index ? io_enq_bits : mem_106; // @[AsyncQueue.scala 47:37]
  assign _GEN_108 = 8'h6b == index ? io_enq_bits : mem_107; // @[AsyncQueue.scala 47:37]
  assign _GEN_109 = 8'h6c == index ? io_enq_bits : mem_108; // @[AsyncQueue.scala 47:37]
  assign _GEN_110 = 8'h6d == index ? io_enq_bits : mem_109; // @[AsyncQueue.scala 47:37]
  assign _GEN_111 = 8'h6e == index ? io_enq_bits : mem_110; // @[AsyncQueue.scala 47:37]
  assign _GEN_112 = 8'h6f == index ? io_enq_bits : mem_111; // @[AsyncQueue.scala 47:37]
  assign _GEN_113 = 8'h70 == index ? io_enq_bits : mem_112; // @[AsyncQueue.scala 47:37]
  assign _GEN_114 = 8'h71 == index ? io_enq_bits : mem_113; // @[AsyncQueue.scala 47:37]
  assign _GEN_115 = 8'h72 == index ? io_enq_bits : mem_114; // @[AsyncQueue.scala 47:37]
  assign _GEN_116 = 8'h73 == index ? io_enq_bits : mem_115; // @[AsyncQueue.scala 47:37]
  assign _GEN_117 = 8'h74 == index ? io_enq_bits : mem_116; // @[AsyncQueue.scala 47:37]
  assign _GEN_118 = 8'h75 == index ? io_enq_bits : mem_117; // @[AsyncQueue.scala 47:37]
  assign _GEN_119 = 8'h76 == index ? io_enq_bits : mem_118; // @[AsyncQueue.scala 47:37]
  assign _GEN_120 = 8'h77 == index ? io_enq_bits : mem_119; // @[AsyncQueue.scala 47:37]
  assign _GEN_121 = 8'h78 == index ? io_enq_bits : mem_120; // @[AsyncQueue.scala 47:37]
  assign _GEN_122 = 8'h79 == index ? io_enq_bits : mem_121; // @[AsyncQueue.scala 47:37]
  assign _GEN_123 = 8'h7a == index ? io_enq_bits : mem_122; // @[AsyncQueue.scala 47:37]
  assign _GEN_124 = 8'h7b == index ? io_enq_bits : mem_123; // @[AsyncQueue.scala 47:37]
  assign _GEN_125 = 8'h7c == index ? io_enq_bits : mem_124; // @[AsyncQueue.scala 47:37]
  assign _GEN_126 = 8'h7d == index ? io_enq_bits : mem_125; // @[AsyncQueue.scala 47:37]
  assign _GEN_127 = 8'h7e == index ? io_enq_bits : mem_126; // @[AsyncQueue.scala 47:37]
  assign _GEN_128 = 8'h7f == index ? io_enq_bits : mem_127; // @[AsyncQueue.scala 47:37]
  assign _GEN_129 = 8'h80 == index ? io_enq_bits : mem_128; // @[AsyncQueue.scala 47:37]
  assign _GEN_130 = 8'h81 == index ? io_enq_bits : mem_129; // @[AsyncQueue.scala 47:37]
  assign _GEN_131 = 8'h82 == index ? io_enq_bits : mem_130; // @[AsyncQueue.scala 47:37]
  assign _GEN_132 = 8'h83 == index ? io_enq_bits : mem_131; // @[AsyncQueue.scala 47:37]
  assign _GEN_133 = 8'h84 == index ? io_enq_bits : mem_132; // @[AsyncQueue.scala 47:37]
  assign _GEN_134 = 8'h85 == index ? io_enq_bits : mem_133; // @[AsyncQueue.scala 47:37]
  assign _GEN_135 = 8'h86 == index ? io_enq_bits : mem_134; // @[AsyncQueue.scala 47:37]
  assign _GEN_136 = 8'h87 == index ? io_enq_bits : mem_135; // @[AsyncQueue.scala 47:37]
  assign _GEN_137 = 8'h88 == index ? io_enq_bits : mem_136; // @[AsyncQueue.scala 47:37]
  assign _GEN_138 = 8'h89 == index ? io_enq_bits : mem_137; // @[AsyncQueue.scala 47:37]
  assign _GEN_139 = 8'h8a == index ? io_enq_bits : mem_138; // @[AsyncQueue.scala 47:37]
  assign _GEN_140 = 8'h8b == index ? io_enq_bits : mem_139; // @[AsyncQueue.scala 47:37]
  assign _GEN_141 = 8'h8c == index ? io_enq_bits : mem_140; // @[AsyncQueue.scala 47:37]
  assign _GEN_142 = 8'h8d == index ? io_enq_bits : mem_141; // @[AsyncQueue.scala 47:37]
  assign _GEN_143 = 8'h8e == index ? io_enq_bits : mem_142; // @[AsyncQueue.scala 47:37]
  assign _GEN_144 = 8'h8f == index ? io_enq_bits : mem_143; // @[AsyncQueue.scala 47:37]
  assign _GEN_145 = 8'h90 == index ? io_enq_bits : mem_144; // @[AsyncQueue.scala 47:37]
  assign _GEN_146 = 8'h91 == index ? io_enq_bits : mem_145; // @[AsyncQueue.scala 47:37]
  assign _GEN_147 = 8'h92 == index ? io_enq_bits : mem_146; // @[AsyncQueue.scala 47:37]
  assign _GEN_148 = 8'h93 == index ? io_enq_bits : mem_147; // @[AsyncQueue.scala 47:37]
  assign _GEN_149 = 8'h94 == index ? io_enq_bits : mem_148; // @[AsyncQueue.scala 47:37]
  assign _GEN_150 = 8'h95 == index ? io_enq_bits : mem_149; // @[AsyncQueue.scala 47:37]
  assign _GEN_151 = 8'h96 == index ? io_enq_bits : mem_150; // @[AsyncQueue.scala 47:37]
  assign _GEN_152 = 8'h97 == index ? io_enq_bits : mem_151; // @[AsyncQueue.scala 47:37]
  assign _GEN_153 = 8'h98 == index ? io_enq_bits : mem_152; // @[AsyncQueue.scala 47:37]
  assign _GEN_154 = 8'h99 == index ? io_enq_bits : mem_153; // @[AsyncQueue.scala 47:37]
  assign _GEN_155 = 8'h9a == index ? io_enq_bits : mem_154; // @[AsyncQueue.scala 47:37]
  assign _GEN_156 = 8'h9b == index ? io_enq_bits : mem_155; // @[AsyncQueue.scala 47:37]
  assign _GEN_157 = 8'h9c == index ? io_enq_bits : mem_156; // @[AsyncQueue.scala 47:37]
  assign _GEN_158 = 8'h9d == index ? io_enq_bits : mem_157; // @[AsyncQueue.scala 47:37]
  assign _GEN_159 = 8'h9e == index ? io_enq_bits : mem_158; // @[AsyncQueue.scala 47:37]
  assign _GEN_160 = 8'h9f == index ? io_enq_bits : mem_159; // @[AsyncQueue.scala 47:37]
  assign _GEN_161 = 8'ha0 == index ? io_enq_bits : mem_160; // @[AsyncQueue.scala 47:37]
  assign _GEN_162 = 8'ha1 == index ? io_enq_bits : mem_161; // @[AsyncQueue.scala 47:37]
  assign _GEN_163 = 8'ha2 == index ? io_enq_bits : mem_162; // @[AsyncQueue.scala 47:37]
  assign _GEN_164 = 8'ha3 == index ? io_enq_bits : mem_163; // @[AsyncQueue.scala 47:37]
  assign _GEN_165 = 8'ha4 == index ? io_enq_bits : mem_164; // @[AsyncQueue.scala 47:37]
  assign _GEN_166 = 8'ha5 == index ? io_enq_bits : mem_165; // @[AsyncQueue.scala 47:37]
  assign _GEN_167 = 8'ha6 == index ? io_enq_bits : mem_166; // @[AsyncQueue.scala 47:37]
  assign _GEN_168 = 8'ha7 == index ? io_enq_bits : mem_167; // @[AsyncQueue.scala 47:37]
  assign _GEN_169 = 8'ha8 == index ? io_enq_bits : mem_168; // @[AsyncQueue.scala 47:37]
  assign _GEN_170 = 8'ha9 == index ? io_enq_bits : mem_169; // @[AsyncQueue.scala 47:37]
  assign _GEN_171 = 8'haa == index ? io_enq_bits : mem_170; // @[AsyncQueue.scala 47:37]
  assign _GEN_172 = 8'hab == index ? io_enq_bits : mem_171; // @[AsyncQueue.scala 47:37]
  assign _GEN_173 = 8'hac == index ? io_enq_bits : mem_172; // @[AsyncQueue.scala 47:37]
  assign _GEN_174 = 8'had == index ? io_enq_bits : mem_173; // @[AsyncQueue.scala 47:37]
  assign _GEN_175 = 8'hae == index ? io_enq_bits : mem_174; // @[AsyncQueue.scala 47:37]
  assign _GEN_176 = 8'haf == index ? io_enq_bits : mem_175; // @[AsyncQueue.scala 47:37]
  assign _GEN_177 = 8'hb0 == index ? io_enq_bits : mem_176; // @[AsyncQueue.scala 47:37]
  assign _GEN_178 = 8'hb1 == index ? io_enq_bits : mem_177; // @[AsyncQueue.scala 47:37]
  assign _GEN_179 = 8'hb2 == index ? io_enq_bits : mem_178; // @[AsyncQueue.scala 47:37]
  assign _GEN_180 = 8'hb3 == index ? io_enq_bits : mem_179; // @[AsyncQueue.scala 47:37]
  assign _GEN_181 = 8'hb4 == index ? io_enq_bits : mem_180; // @[AsyncQueue.scala 47:37]
  assign _GEN_182 = 8'hb5 == index ? io_enq_bits : mem_181; // @[AsyncQueue.scala 47:37]
  assign _GEN_183 = 8'hb6 == index ? io_enq_bits : mem_182; // @[AsyncQueue.scala 47:37]
  assign _GEN_184 = 8'hb7 == index ? io_enq_bits : mem_183; // @[AsyncQueue.scala 47:37]
  assign _GEN_185 = 8'hb8 == index ? io_enq_bits : mem_184; // @[AsyncQueue.scala 47:37]
  assign _GEN_186 = 8'hb9 == index ? io_enq_bits : mem_185; // @[AsyncQueue.scala 47:37]
  assign _GEN_187 = 8'hba == index ? io_enq_bits : mem_186; // @[AsyncQueue.scala 47:37]
  assign _GEN_188 = 8'hbb == index ? io_enq_bits : mem_187; // @[AsyncQueue.scala 47:37]
  assign _GEN_189 = 8'hbc == index ? io_enq_bits : mem_188; // @[AsyncQueue.scala 47:37]
  assign _GEN_190 = 8'hbd == index ? io_enq_bits : mem_189; // @[AsyncQueue.scala 47:37]
  assign _GEN_191 = 8'hbe == index ? io_enq_bits : mem_190; // @[AsyncQueue.scala 47:37]
  assign _GEN_192 = 8'hbf == index ? io_enq_bits : mem_191; // @[AsyncQueue.scala 47:37]
  assign _GEN_193 = 8'hc0 == index ? io_enq_bits : mem_192; // @[AsyncQueue.scala 47:37]
  assign _GEN_194 = 8'hc1 == index ? io_enq_bits : mem_193; // @[AsyncQueue.scala 47:37]
  assign _GEN_195 = 8'hc2 == index ? io_enq_bits : mem_194; // @[AsyncQueue.scala 47:37]
  assign _GEN_196 = 8'hc3 == index ? io_enq_bits : mem_195; // @[AsyncQueue.scala 47:37]
  assign _GEN_197 = 8'hc4 == index ? io_enq_bits : mem_196; // @[AsyncQueue.scala 47:37]
  assign _GEN_198 = 8'hc5 == index ? io_enq_bits : mem_197; // @[AsyncQueue.scala 47:37]
  assign _GEN_199 = 8'hc6 == index ? io_enq_bits : mem_198; // @[AsyncQueue.scala 47:37]
  assign _GEN_200 = 8'hc7 == index ? io_enq_bits : mem_199; // @[AsyncQueue.scala 47:37]
  assign _GEN_201 = 8'hc8 == index ? io_enq_bits : mem_200; // @[AsyncQueue.scala 47:37]
  assign _GEN_202 = 8'hc9 == index ? io_enq_bits : mem_201; // @[AsyncQueue.scala 47:37]
  assign _GEN_203 = 8'hca == index ? io_enq_bits : mem_202; // @[AsyncQueue.scala 47:37]
  assign _GEN_204 = 8'hcb == index ? io_enq_bits : mem_203; // @[AsyncQueue.scala 47:37]
  assign _GEN_205 = 8'hcc == index ? io_enq_bits : mem_204; // @[AsyncQueue.scala 47:37]
  assign _GEN_206 = 8'hcd == index ? io_enq_bits : mem_205; // @[AsyncQueue.scala 47:37]
  assign _GEN_207 = 8'hce == index ? io_enq_bits : mem_206; // @[AsyncQueue.scala 47:37]
  assign _GEN_208 = 8'hcf == index ? io_enq_bits : mem_207; // @[AsyncQueue.scala 47:37]
  assign _GEN_209 = 8'hd0 == index ? io_enq_bits : mem_208; // @[AsyncQueue.scala 47:37]
  assign _GEN_210 = 8'hd1 == index ? io_enq_bits : mem_209; // @[AsyncQueue.scala 47:37]
  assign _GEN_211 = 8'hd2 == index ? io_enq_bits : mem_210; // @[AsyncQueue.scala 47:37]
  assign _GEN_212 = 8'hd3 == index ? io_enq_bits : mem_211; // @[AsyncQueue.scala 47:37]
  assign _GEN_213 = 8'hd4 == index ? io_enq_bits : mem_212; // @[AsyncQueue.scala 47:37]
  assign _GEN_214 = 8'hd5 == index ? io_enq_bits : mem_213; // @[AsyncQueue.scala 47:37]
  assign _GEN_215 = 8'hd6 == index ? io_enq_bits : mem_214; // @[AsyncQueue.scala 47:37]
  assign _GEN_216 = 8'hd7 == index ? io_enq_bits : mem_215; // @[AsyncQueue.scala 47:37]
  assign _GEN_217 = 8'hd8 == index ? io_enq_bits : mem_216; // @[AsyncQueue.scala 47:37]
  assign _GEN_218 = 8'hd9 == index ? io_enq_bits : mem_217; // @[AsyncQueue.scala 47:37]
  assign _GEN_219 = 8'hda == index ? io_enq_bits : mem_218; // @[AsyncQueue.scala 47:37]
  assign _GEN_220 = 8'hdb == index ? io_enq_bits : mem_219; // @[AsyncQueue.scala 47:37]
  assign _GEN_221 = 8'hdc == index ? io_enq_bits : mem_220; // @[AsyncQueue.scala 47:37]
  assign _GEN_222 = 8'hdd == index ? io_enq_bits : mem_221; // @[AsyncQueue.scala 47:37]
  assign _GEN_223 = 8'hde == index ? io_enq_bits : mem_222; // @[AsyncQueue.scala 47:37]
  assign _GEN_224 = 8'hdf == index ? io_enq_bits : mem_223; // @[AsyncQueue.scala 47:37]
  assign _GEN_225 = 8'he0 == index ? io_enq_bits : mem_224; // @[AsyncQueue.scala 47:37]
  assign _GEN_226 = 8'he1 == index ? io_enq_bits : mem_225; // @[AsyncQueue.scala 47:37]
  assign _GEN_227 = 8'he2 == index ? io_enq_bits : mem_226; // @[AsyncQueue.scala 47:37]
  assign _GEN_228 = 8'he3 == index ? io_enq_bits : mem_227; // @[AsyncQueue.scala 47:37]
  assign _GEN_229 = 8'he4 == index ? io_enq_bits : mem_228; // @[AsyncQueue.scala 47:37]
  assign _GEN_230 = 8'he5 == index ? io_enq_bits : mem_229; // @[AsyncQueue.scala 47:37]
  assign _GEN_231 = 8'he6 == index ? io_enq_bits : mem_230; // @[AsyncQueue.scala 47:37]
  assign _GEN_232 = 8'he7 == index ? io_enq_bits : mem_231; // @[AsyncQueue.scala 47:37]
  assign _GEN_233 = 8'he8 == index ? io_enq_bits : mem_232; // @[AsyncQueue.scala 47:37]
  assign _GEN_234 = 8'he9 == index ? io_enq_bits : mem_233; // @[AsyncQueue.scala 47:37]
  assign _GEN_235 = 8'hea == index ? io_enq_bits : mem_234; // @[AsyncQueue.scala 47:37]
  assign _GEN_236 = 8'heb == index ? io_enq_bits : mem_235; // @[AsyncQueue.scala 47:37]
  assign _GEN_237 = 8'hec == index ? io_enq_bits : mem_236; // @[AsyncQueue.scala 47:37]
  assign _GEN_238 = 8'hed == index ? io_enq_bits : mem_237; // @[AsyncQueue.scala 47:37]
  assign _GEN_239 = 8'hee == index ? io_enq_bits : mem_238; // @[AsyncQueue.scala 47:37]
  assign _GEN_240 = 8'hef == index ? io_enq_bits : mem_239; // @[AsyncQueue.scala 47:37]
  assign _GEN_241 = 8'hf0 == index ? io_enq_bits : mem_240; // @[AsyncQueue.scala 47:37]
  assign _GEN_242 = 8'hf1 == index ? io_enq_bits : mem_241; // @[AsyncQueue.scala 47:37]
  assign _GEN_243 = 8'hf2 == index ? io_enq_bits : mem_242; // @[AsyncQueue.scala 47:37]
  assign _GEN_244 = 8'hf3 == index ? io_enq_bits : mem_243; // @[AsyncQueue.scala 47:37]
  assign _GEN_245 = 8'hf4 == index ? io_enq_bits : mem_244; // @[AsyncQueue.scala 47:37]
  assign _GEN_246 = 8'hf5 == index ? io_enq_bits : mem_245; // @[AsyncQueue.scala 47:37]
  assign _GEN_247 = 8'hf6 == index ? io_enq_bits : mem_246; // @[AsyncQueue.scala 47:37]
  assign _GEN_248 = 8'hf7 == index ? io_enq_bits : mem_247; // @[AsyncQueue.scala 47:37]
  assign _GEN_249 = 8'hf8 == index ? io_enq_bits : mem_248; // @[AsyncQueue.scala 47:37]
  assign _GEN_250 = 8'hf9 == index ? io_enq_bits : mem_249; // @[AsyncQueue.scala 47:37]
  assign _GEN_251 = 8'hfa == index ? io_enq_bits : mem_250; // @[AsyncQueue.scala 47:37]
  assign _GEN_252 = 8'hfb == index ? io_enq_bits : mem_251; // @[AsyncQueue.scala 47:37]
  assign _GEN_253 = 8'hfc == index ? io_enq_bits : mem_252; // @[AsyncQueue.scala 47:37]
  assign _GEN_254 = 8'hfd == index ? io_enq_bits : mem_253; // @[AsyncQueue.scala 47:37]
  assign _GEN_255 = 8'hfe == index ? io_enq_bits : mem_254; // @[AsyncQueue.scala 47:37]
  assign _GEN_256 = 8'hff == index ? io_enq_bits : mem_255; // @[AsyncQueue.scala 47:37]
  assign _GEN_257 = _T_536 ? _GEN_1 : mem_0; // @[AsyncQueue.scala 47:24]
  assign _GEN_258 = _T_536 ? _GEN_2 : mem_1; // @[AsyncQueue.scala 47:24]
  assign _GEN_259 = _T_536 ? _GEN_3 : mem_2; // @[AsyncQueue.scala 47:24]
  assign _GEN_260 = _T_536 ? _GEN_4 : mem_3; // @[AsyncQueue.scala 47:24]
  assign _GEN_261 = _T_536 ? _GEN_5 : mem_4; // @[AsyncQueue.scala 47:24]
  assign _GEN_262 = _T_536 ? _GEN_6 : mem_5; // @[AsyncQueue.scala 47:24]
  assign _GEN_263 = _T_536 ? _GEN_7 : mem_6; // @[AsyncQueue.scala 47:24]
  assign _GEN_264 = _T_536 ? _GEN_8 : mem_7; // @[AsyncQueue.scala 47:24]
  assign _GEN_265 = _T_536 ? _GEN_9 : mem_8; // @[AsyncQueue.scala 47:24]
  assign _GEN_266 = _T_536 ? _GEN_10 : mem_9; // @[AsyncQueue.scala 47:24]
  assign _GEN_267 = _T_536 ? _GEN_11 : mem_10; // @[AsyncQueue.scala 47:24]
  assign _GEN_268 = _T_536 ? _GEN_12 : mem_11; // @[AsyncQueue.scala 47:24]
  assign _GEN_269 = _T_536 ? _GEN_13 : mem_12; // @[AsyncQueue.scala 47:24]
  assign _GEN_270 = _T_536 ? _GEN_14 : mem_13; // @[AsyncQueue.scala 47:24]
  assign _GEN_271 = _T_536 ? _GEN_15 : mem_14; // @[AsyncQueue.scala 47:24]
  assign _GEN_272 = _T_536 ? _GEN_16 : mem_15; // @[AsyncQueue.scala 47:24]
  assign _GEN_273 = _T_536 ? _GEN_17 : mem_16; // @[AsyncQueue.scala 47:24]
  assign _GEN_274 = _T_536 ? _GEN_18 : mem_17; // @[AsyncQueue.scala 47:24]
  assign _GEN_275 = _T_536 ? _GEN_19 : mem_18; // @[AsyncQueue.scala 47:24]
  assign _GEN_276 = _T_536 ? _GEN_20 : mem_19; // @[AsyncQueue.scala 47:24]
  assign _GEN_277 = _T_536 ? _GEN_21 : mem_20; // @[AsyncQueue.scala 47:24]
  assign _GEN_278 = _T_536 ? _GEN_22 : mem_21; // @[AsyncQueue.scala 47:24]
  assign _GEN_279 = _T_536 ? _GEN_23 : mem_22; // @[AsyncQueue.scala 47:24]
  assign _GEN_280 = _T_536 ? _GEN_24 : mem_23; // @[AsyncQueue.scala 47:24]
  assign _GEN_281 = _T_536 ? _GEN_25 : mem_24; // @[AsyncQueue.scala 47:24]
  assign _GEN_282 = _T_536 ? _GEN_26 : mem_25; // @[AsyncQueue.scala 47:24]
  assign _GEN_283 = _T_536 ? _GEN_27 : mem_26; // @[AsyncQueue.scala 47:24]
  assign _GEN_284 = _T_536 ? _GEN_28 : mem_27; // @[AsyncQueue.scala 47:24]
  assign _GEN_285 = _T_536 ? _GEN_29 : mem_28; // @[AsyncQueue.scala 47:24]
  assign _GEN_286 = _T_536 ? _GEN_30 : mem_29; // @[AsyncQueue.scala 47:24]
  assign _GEN_287 = _T_536 ? _GEN_31 : mem_30; // @[AsyncQueue.scala 47:24]
  assign _GEN_288 = _T_536 ? _GEN_32 : mem_31; // @[AsyncQueue.scala 47:24]
  assign _GEN_289 = _T_536 ? _GEN_33 : mem_32; // @[AsyncQueue.scala 47:24]
  assign _GEN_290 = _T_536 ? _GEN_34 : mem_33; // @[AsyncQueue.scala 47:24]
  assign _GEN_291 = _T_536 ? _GEN_35 : mem_34; // @[AsyncQueue.scala 47:24]
  assign _GEN_292 = _T_536 ? _GEN_36 : mem_35; // @[AsyncQueue.scala 47:24]
  assign _GEN_293 = _T_536 ? _GEN_37 : mem_36; // @[AsyncQueue.scala 47:24]
  assign _GEN_294 = _T_536 ? _GEN_38 : mem_37; // @[AsyncQueue.scala 47:24]
  assign _GEN_295 = _T_536 ? _GEN_39 : mem_38; // @[AsyncQueue.scala 47:24]
  assign _GEN_296 = _T_536 ? _GEN_40 : mem_39; // @[AsyncQueue.scala 47:24]
  assign _GEN_297 = _T_536 ? _GEN_41 : mem_40; // @[AsyncQueue.scala 47:24]
  assign _GEN_298 = _T_536 ? _GEN_42 : mem_41; // @[AsyncQueue.scala 47:24]
  assign _GEN_299 = _T_536 ? _GEN_43 : mem_42; // @[AsyncQueue.scala 47:24]
  assign _GEN_300 = _T_536 ? _GEN_44 : mem_43; // @[AsyncQueue.scala 47:24]
  assign _GEN_301 = _T_536 ? _GEN_45 : mem_44; // @[AsyncQueue.scala 47:24]
  assign _GEN_302 = _T_536 ? _GEN_46 : mem_45; // @[AsyncQueue.scala 47:24]
  assign _GEN_303 = _T_536 ? _GEN_47 : mem_46; // @[AsyncQueue.scala 47:24]
  assign _GEN_304 = _T_536 ? _GEN_48 : mem_47; // @[AsyncQueue.scala 47:24]
  assign _GEN_305 = _T_536 ? _GEN_49 : mem_48; // @[AsyncQueue.scala 47:24]
  assign _GEN_306 = _T_536 ? _GEN_50 : mem_49; // @[AsyncQueue.scala 47:24]
  assign _GEN_307 = _T_536 ? _GEN_51 : mem_50; // @[AsyncQueue.scala 47:24]
  assign _GEN_308 = _T_536 ? _GEN_52 : mem_51; // @[AsyncQueue.scala 47:24]
  assign _GEN_309 = _T_536 ? _GEN_53 : mem_52; // @[AsyncQueue.scala 47:24]
  assign _GEN_310 = _T_536 ? _GEN_54 : mem_53; // @[AsyncQueue.scala 47:24]
  assign _GEN_311 = _T_536 ? _GEN_55 : mem_54; // @[AsyncQueue.scala 47:24]
  assign _GEN_312 = _T_536 ? _GEN_56 : mem_55; // @[AsyncQueue.scala 47:24]
  assign _GEN_313 = _T_536 ? _GEN_57 : mem_56; // @[AsyncQueue.scala 47:24]
  assign _GEN_314 = _T_536 ? _GEN_58 : mem_57; // @[AsyncQueue.scala 47:24]
  assign _GEN_315 = _T_536 ? _GEN_59 : mem_58; // @[AsyncQueue.scala 47:24]
  assign _GEN_316 = _T_536 ? _GEN_60 : mem_59; // @[AsyncQueue.scala 47:24]
  assign _GEN_317 = _T_536 ? _GEN_61 : mem_60; // @[AsyncQueue.scala 47:24]
  assign _GEN_318 = _T_536 ? _GEN_62 : mem_61; // @[AsyncQueue.scala 47:24]
  assign _GEN_319 = _T_536 ? _GEN_63 : mem_62; // @[AsyncQueue.scala 47:24]
  assign _GEN_320 = _T_536 ? _GEN_64 : mem_63; // @[AsyncQueue.scala 47:24]
  assign _GEN_321 = _T_536 ? _GEN_65 : mem_64; // @[AsyncQueue.scala 47:24]
  assign _GEN_322 = _T_536 ? _GEN_66 : mem_65; // @[AsyncQueue.scala 47:24]
  assign _GEN_323 = _T_536 ? _GEN_67 : mem_66; // @[AsyncQueue.scala 47:24]
  assign _GEN_324 = _T_536 ? _GEN_68 : mem_67; // @[AsyncQueue.scala 47:24]
  assign _GEN_325 = _T_536 ? _GEN_69 : mem_68; // @[AsyncQueue.scala 47:24]
  assign _GEN_326 = _T_536 ? _GEN_70 : mem_69; // @[AsyncQueue.scala 47:24]
  assign _GEN_327 = _T_536 ? _GEN_71 : mem_70; // @[AsyncQueue.scala 47:24]
  assign _GEN_328 = _T_536 ? _GEN_72 : mem_71; // @[AsyncQueue.scala 47:24]
  assign _GEN_329 = _T_536 ? _GEN_73 : mem_72; // @[AsyncQueue.scala 47:24]
  assign _GEN_330 = _T_536 ? _GEN_74 : mem_73; // @[AsyncQueue.scala 47:24]
  assign _GEN_331 = _T_536 ? _GEN_75 : mem_74; // @[AsyncQueue.scala 47:24]
  assign _GEN_332 = _T_536 ? _GEN_76 : mem_75; // @[AsyncQueue.scala 47:24]
  assign _GEN_333 = _T_536 ? _GEN_77 : mem_76; // @[AsyncQueue.scala 47:24]
  assign _GEN_334 = _T_536 ? _GEN_78 : mem_77; // @[AsyncQueue.scala 47:24]
  assign _GEN_335 = _T_536 ? _GEN_79 : mem_78; // @[AsyncQueue.scala 47:24]
  assign _GEN_336 = _T_536 ? _GEN_80 : mem_79; // @[AsyncQueue.scala 47:24]
  assign _GEN_337 = _T_536 ? _GEN_81 : mem_80; // @[AsyncQueue.scala 47:24]
  assign _GEN_338 = _T_536 ? _GEN_82 : mem_81; // @[AsyncQueue.scala 47:24]
  assign _GEN_339 = _T_536 ? _GEN_83 : mem_82; // @[AsyncQueue.scala 47:24]
  assign _GEN_340 = _T_536 ? _GEN_84 : mem_83; // @[AsyncQueue.scala 47:24]
  assign _GEN_341 = _T_536 ? _GEN_85 : mem_84; // @[AsyncQueue.scala 47:24]
  assign _GEN_342 = _T_536 ? _GEN_86 : mem_85; // @[AsyncQueue.scala 47:24]
  assign _GEN_343 = _T_536 ? _GEN_87 : mem_86; // @[AsyncQueue.scala 47:24]
  assign _GEN_344 = _T_536 ? _GEN_88 : mem_87; // @[AsyncQueue.scala 47:24]
  assign _GEN_345 = _T_536 ? _GEN_89 : mem_88; // @[AsyncQueue.scala 47:24]
  assign _GEN_346 = _T_536 ? _GEN_90 : mem_89; // @[AsyncQueue.scala 47:24]
  assign _GEN_347 = _T_536 ? _GEN_91 : mem_90; // @[AsyncQueue.scala 47:24]
  assign _GEN_348 = _T_536 ? _GEN_92 : mem_91; // @[AsyncQueue.scala 47:24]
  assign _GEN_349 = _T_536 ? _GEN_93 : mem_92; // @[AsyncQueue.scala 47:24]
  assign _GEN_350 = _T_536 ? _GEN_94 : mem_93; // @[AsyncQueue.scala 47:24]
  assign _GEN_351 = _T_536 ? _GEN_95 : mem_94; // @[AsyncQueue.scala 47:24]
  assign _GEN_352 = _T_536 ? _GEN_96 : mem_95; // @[AsyncQueue.scala 47:24]
  assign _GEN_353 = _T_536 ? _GEN_97 : mem_96; // @[AsyncQueue.scala 47:24]
  assign _GEN_354 = _T_536 ? _GEN_98 : mem_97; // @[AsyncQueue.scala 47:24]
  assign _GEN_355 = _T_536 ? _GEN_99 : mem_98; // @[AsyncQueue.scala 47:24]
  assign _GEN_356 = _T_536 ? _GEN_100 : mem_99; // @[AsyncQueue.scala 47:24]
  assign _GEN_357 = _T_536 ? _GEN_101 : mem_100; // @[AsyncQueue.scala 47:24]
  assign _GEN_358 = _T_536 ? _GEN_102 : mem_101; // @[AsyncQueue.scala 47:24]
  assign _GEN_359 = _T_536 ? _GEN_103 : mem_102; // @[AsyncQueue.scala 47:24]
  assign _GEN_360 = _T_536 ? _GEN_104 : mem_103; // @[AsyncQueue.scala 47:24]
  assign _GEN_361 = _T_536 ? _GEN_105 : mem_104; // @[AsyncQueue.scala 47:24]
  assign _GEN_362 = _T_536 ? _GEN_106 : mem_105; // @[AsyncQueue.scala 47:24]
  assign _GEN_363 = _T_536 ? _GEN_107 : mem_106; // @[AsyncQueue.scala 47:24]
  assign _GEN_364 = _T_536 ? _GEN_108 : mem_107; // @[AsyncQueue.scala 47:24]
  assign _GEN_365 = _T_536 ? _GEN_109 : mem_108; // @[AsyncQueue.scala 47:24]
  assign _GEN_366 = _T_536 ? _GEN_110 : mem_109; // @[AsyncQueue.scala 47:24]
  assign _GEN_367 = _T_536 ? _GEN_111 : mem_110; // @[AsyncQueue.scala 47:24]
  assign _GEN_368 = _T_536 ? _GEN_112 : mem_111; // @[AsyncQueue.scala 47:24]
  assign _GEN_369 = _T_536 ? _GEN_113 : mem_112; // @[AsyncQueue.scala 47:24]
  assign _GEN_370 = _T_536 ? _GEN_114 : mem_113; // @[AsyncQueue.scala 47:24]
  assign _GEN_371 = _T_536 ? _GEN_115 : mem_114; // @[AsyncQueue.scala 47:24]
  assign _GEN_372 = _T_536 ? _GEN_116 : mem_115; // @[AsyncQueue.scala 47:24]
  assign _GEN_373 = _T_536 ? _GEN_117 : mem_116; // @[AsyncQueue.scala 47:24]
  assign _GEN_374 = _T_536 ? _GEN_118 : mem_117; // @[AsyncQueue.scala 47:24]
  assign _GEN_375 = _T_536 ? _GEN_119 : mem_118; // @[AsyncQueue.scala 47:24]
  assign _GEN_376 = _T_536 ? _GEN_120 : mem_119; // @[AsyncQueue.scala 47:24]
  assign _GEN_377 = _T_536 ? _GEN_121 : mem_120; // @[AsyncQueue.scala 47:24]
  assign _GEN_378 = _T_536 ? _GEN_122 : mem_121; // @[AsyncQueue.scala 47:24]
  assign _GEN_379 = _T_536 ? _GEN_123 : mem_122; // @[AsyncQueue.scala 47:24]
  assign _GEN_380 = _T_536 ? _GEN_124 : mem_123; // @[AsyncQueue.scala 47:24]
  assign _GEN_381 = _T_536 ? _GEN_125 : mem_124; // @[AsyncQueue.scala 47:24]
  assign _GEN_382 = _T_536 ? _GEN_126 : mem_125; // @[AsyncQueue.scala 47:24]
  assign _GEN_383 = _T_536 ? _GEN_127 : mem_126; // @[AsyncQueue.scala 47:24]
  assign _GEN_384 = _T_536 ? _GEN_128 : mem_127; // @[AsyncQueue.scala 47:24]
  assign _GEN_385 = _T_536 ? _GEN_129 : mem_128; // @[AsyncQueue.scala 47:24]
  assign _GEN_386 = _T_536 ? _GEN_130 : mem_129; // @[AsyncQueue.scala 47:24]
  assign _GEN_387 = _T_536 ? _GEN_131 : mem_130; // @[AsyncQueue.scala 47:24]
  assign _GEN_388 = _T_536 ? _GEN_132 : mem_131; // @[AsyncQueue.scala 47:24]
  assign _GEN_389 = _T_536 ? _GEN_133 : mem_132; // @[AsyncQueue.scala 47:24]
  assign _GEN_390 = _T_536 ? _GEN_134 : mem_133; // @[AsyncQueue.scala 47:24]
  assign _GEN_391 = _T_536 ? _GEN_135 : mem_134; // @[AsyncQueue.scala 47:24]
  assign _GEN_392 = _T_536 ? _GEN_136 : mem_135; // @[AsyncQueue.scala 47:24]
  assign _GEN_393 = _T_536 ? _GEN_137 : mem_136; // @[AsyncQueue.scala 47:24]
  assign _GEN_394 = _T_536 ? _GEN_138 : mem_137; // @[AsyncQueue.scala 47:24]
  assign _GEN_395 = _T_536 ? _GEN_139 : mem_138; // @[AsyncQueue.scala 47:24]
  assign _GEN_396 = _T_536 ? _GEN_140 : mem_139; // @[AsyncQueue.scala 47:24]
  assign _GEN_397 = _T_536 ? _GEN_141 : mem_140; // @[AsyncQueue.scala 47:24]
  assign _GEN_398 = _T_536 ? _GEN_142 : mem_141; // @[AsyncQueue.scala 47:24]
  assign _GEN_399 = _T_536 ? _GEN_143 : mem_142; // @[AsyncQueue.scala 47:24]
  assign _GEN_400 = _T_536 ? _GEN_144 : mem_143; // @[AsyncQueue.scala 47:24]
  assign _GEN_401 = _T_536 ? _GEN_145 : mem_144; // @[AsyncQueue.scala 47:24]
  assign _GEN_402 = _T_536 ? _GEN_146 : mem_145; // @[AsyncQueue.scala 47:24]
  assign _GEN_403 = _T_536 ? _GEN_147 : mem_146; // @[AsyncQueue.scala 47:24]
  assign _GEN_404 = _T_536 ? _GEN_148 : mem_147; // @[AsyncQueue.scala 47:24]
  assign _GEN_405 = _T_536 ? _GEN_149 : mem_148; // @[AsyncQueue.scala 47:24]
  assign _GEN_406 = _T_536 ? _GEN_150 : mem_149; // @[AsyncQueue.scala 47:24]
  assign _GEN_407 = _T_536 ? _GEN_151 : mem_150; // @[AsyncQueue.scala 47:24]
  assign _GEN_408 = _T_536 ? _GEN_152 : mem_151; // @[AsyncQueue.scala 47:24]
  assign _GEN_409 = _T_536 ? _GEN_153 : mem_152; // @[AsyncQueue.scala 47:24]
  assign _GEN_410 = _T_536 ? _GEN_154 : mem_153; // @[AsyncQueue.scala 47:24]
  assign _GEN_411 = _T_536 ? _GEN_155 : mem_154; // @[AsyncQueue.scala 47:24]
  assign _GEN_412 = _T_536 ? _GEN_156 : mem_155; // @[AsyncQueue.scala 47:24]
  assign _GEN_413 = _T_536 ? _GEN_157 : mem_156; // @[AsyncQueue.scala 47:24]
  assign _GEN_414 = _T_536 ? _GEN_158 : mem_157; // @[AsyncQueue.scala 47:24]
  assign _GEN_415 = _T_536 ? _GEN_159 : mem_158; // @[AsyncQueue.scala 47:24]
  assign _GEN_416 = _T_536 ? _GEN_160 : mem_159; // @[AsyncQueue.scala 47:24]
  assign _GEN_417 = _T_536 ? _GEN_161 : mem_160; // @[AsyncQueue.scala 47:24]
  assign _GEN_418 = _T_536 ? _GEN_162 : mem_161; // @[AsyncQueue.scala 47:24]
  assign _GEN_419 = _T_536 ? _GEN_163 : mem_162; // @[AsyncQueue.scala 47:24]
  assign _GEN_420 = _T_536 ? _GEN_164 : mem_163; // @[AsyncQueue.scala 47:24]
  assign _GEN_421 = _T_536 ? _GEN_165 : mem_164; // @[AsyncQueue.scala 47:24]
  assign _GEN_422 = _T_536 ? _GEN_166 : mem_165; // @[AsyncQueue.scala 47:24]
  assign _GEN_423 = _T_536 ? _GEN_167 : mem_166; // @[AsyncQueue.scala 47:24]
  assign _GEN_424 = _T_536 ? _GEN_168 : mem_167; // @[AsyncQueue.scala 47:24]
  assign _GEN_425 = _T_536 ? _GEN_169 : mem_168; // @[AsyncQueue.scala 47:24]
  assign _GEN_426 = _T_536 ? _GEN_170 : mem_169; // @[AsyncQueue.scala 47:24]
  assign _GEN_427 = _T_536 ? _GEN_171 : mem_170; // @[AsyncQueue.scala 47:24]
  assign _GEN_428 = _T_536 ? _GEN_172 : mem_171; // @[AsyncQueue.scala 47:24]
  assign _GEN_429 = _T_536 ? _GEN_173 : mem_172; // @[AsyncQueue.scala 47:24]
  assign _GEN_430 = _T_536 ? _GEN_174 : mem_173; // @[AsyncQueue.scala 47:24]
  assign _GEN_431 = _T_536 ? _GEN_175 : mem_174; // @[AsyncQueue.scala 47:24]
  assign _GEN_432 = _T_536 ? _GEN_176 : mem_175; // @[AsyncQueue.scala 47:24]
  assign _GEN_433 = _T_536 ? _GEN_177 : mem_176; // @[AsyncQueue.scala 47:24]
  assign _GEN_434 = _T_536 ? _GEN_178 : mem_177; // @[AsyncQueue.scala 47:24]
  assign _GEN_435 = _T_536 ? _GEN_179 : mem_178; // @[AsyncQueue.scala 47:24]
  assign _GEN_436 = _T_536 ? _GEN_180 : mem_179; // @[AsyncQueue.scala 47:24]
  assign _GEN_437 = _T_536 ? _GEN_181 : mem_180; // @[AsyncQueue.scala 47:24]
  assign _GEN_438 = _T_536 ? _GEN_182 : mem_181; // @[AsyncQueue.scala 47:24]
  assign _GEN_439 = _T_536 ? _GEN_183 : mem_182; // @[AsyncQueue.scala 47:24]
  assign _GEN_440 = _T_536 ? _GEN_184 : mem_183; // @[AsyncQueue.scala 47:24]
  assign _GEN_441 = _T_536 ? _GEN_185 : mem_184; // @[AsyncQueue.scala 47:24]
  assign _GEN_442 = _T_536 ? _GEN_186 : mem_185; // @[AsyncQueue.scala 47:24]
  assign _GEN_443 = _T_536 ? _GEN_187 : mem_186; // @[AsyncQueue.scala 47:24]
  assign _GEN_444 = _T_536 ? _GEN_188 : mem_187; // @[AsyncQueue.scala 47:24]
  assign _GEN_445 = _T_536 ? _GEN_189 : mem_188; // @[AsyncQueue.scala 47:24]
  assign _GEN_446 = _T_536 ? _GEN_190 : mem_189; // @[AsyncQueue.scala 47:24]
  assign _GEN_447 = _T_536 ? _GEN_191 : mem_190; // @[AsyncQueue.scala 47:24]
  assign _GEN_448 = _T_536 ? _GEN_192 : mem_191; // @[AsyncQueue.scala 47:24]
  assign _GEN_449 = _T_536 ? _GEN_193 : mem_192; // @[AsyncQueue.scala 47:24]
  assign _GEN_450 = _T_536 ? _GEN_194 : mem_193; // @[AsyncQueue.scala 47:24]
  assign _GEN_451 = _T_536 ? _GEN_195 : mem_194; // @[AsyncQueue.scala 47:24]
  assign _GEN_452 = _T_536 ? _GEN_196 : mem_195; // @[AsyncQueue.scala 47:24]
  assign _GEN_453 = _T_536 ? _GEN_197 : mem_196; // @[AsyncQueue.scala 47:24]
  assign _GEN_454 = _T_536 ? _GEN_198 : mem_197; // @[AsyncQueue.scala 47:24]
  assign _GEN_455 = _T_536 ? _GEN_199 : mem_198; // @[AsyncQueue.scala 47:24]
  assign _GEN_456 = _T_536 ? _GEN_200 : mem_199; // @[AsyncQueue.scala 47:24]
  assign _GEN_457 = _T_536 ? _GEN_201 : mem_200; // @[AsyncQueue.scala 47:24]
  assign _GEN_458 = _T_536 ? _GEN_202 : mem_201; // @[AsyncQueue.scala 47:24]
  assign _GEN_459 = _T_536 ? _GEN_203 : mem_202; // @[AsyncQueue.scala 47:24]
  assign _GEN_460 = _T_536 ? _GEN_204 : mem_203; // @[AsyncQueue.scala 47:24]
  assign _GEN_461 = _T_536 ? _GEN_205 : mem_204; // @[AsyncQueue.scala 47:24]
  assign _GEN_462 = _T_536 ? _GEN_206 : mem_205; // @[AsyncQueue.scala 47:24]
  assign _GEN_463 = _T_536 ? _GEN_207 : mem_206; // @[AsyncQueue.scala 47:24]
  assign _GEN_464 = _T_536 ? _GEN_208 : mem_207; // @[AsyncQueue.scala 47:24]
  assign _GEN_465 = _T_536 ? _GEN_209 : mem_208; // @[AsyncQueue.scala 47:24]
  assign _GEN_466 = _T_536 ? _GEN_210 : mem_209; // @[AsyncQueue.scala 47:24]
  assign _GEN_467 = _T_536 ? _GEN_211 : mem_210; // @[AsyncQueue.scala 47:24]
  assign _GEN_468 = _T_536 ? _GEN_212 : mem_211; // @[AsyncQueue.scala 47:24]
  assign _GEN_469 = _T_536 ? _GEN_213 : mem_212; // @[AsyncQueue.scala 47:24]
  assign _GEN_470 = _T_536 ? _GEN_214 : mem_213; // @[AsyncQueue.scala 47:24]
  assign _GEN_471 = _T_536 ? _GEN_215 : mem_214; // @[AsyncQueue.scala 47:24]
  assign _GEN_472 = _T_536 ? _GEN_216 : mem_215; // @[AsyncQueue.scala 47:24]
  assign _GEN_473 = _T_536 ? _GEN_217 : mem_216; // @[AsyncQueue.scala 47:24]
  assign _GEN_474 = _T_536 ? _GEN_218 : mem_217; // @[AsyncQueue.scala 47:24]
  assign _GEN_475 = _T_536 ? _GEN_219 : mem_218; // @[AsyncQueue.scala 47:24]
  assign _GEN_476 = _T_536 ? _GEN_220 : mem_219; // @[AsyncQueue.scala 47:24]
  assign _GEN_477 = _T_536 ? _GEN_221 : mem_220; // @[AsyncQueue.scala 47:24]
  assign _GEN_478 = _T_536 ? _GEN_222 : mem_221; // @[AsyncQueue.scala 47:24]
  assign _GEN_479 = _T_536 ? _GEN_223 : mem_222; // @[AsyncQueue.scala 47:24]
  assign _GEN_480 = _T_536 ? _GEN_224 : mem_223; // @[AsyncQueue.scala 47:24]
  assign _GEN_481 = _T_536 ? _GEN_225 : mem_224; // @[AsyncQueue.scala 47:24]
  assign _GEN_482 = _T_536 ? _GEN_226 : mem_225; // @[AsyncQueue.scala 47:24]
  assign _GEN_483 = _T_536 ? _GEN_227 : mem_226; // @[AsyncQueue.scala 47:24]
  assign _GEN_484 = _T_536 ? _GEN_228 : mem_227; // @[AsyncQueue.scala 47:24]
  assign _GEN_485 = _T_536 ? _GEN_229 : mem_228; // @[AsyncQueue.scala 47:24]
  assign _GEN_486 = _T_536 ? _GEN_230 : mem_229; // @[AsyncQueue.scala 47:24]
  assign _GEN_487 = _T_536 ? _GEN_231 : mem_230; // @[AsyncQueue.scala 47:24]
  assign _GEN_488 = _T_536 ? _GEN_232 : mem_231; // @[AsyncQueue.scala 47:24]
  assign _GEN_489 = _T_536 ? _GEN_233 : mem_232; // @[AsyncQueue.scala 47:24]
  assign _GEN_490 = _T_536 ? _GEN_234 : mem_233; // @[AsyncQueue.scala 47:24]
  assign _GEN_491 = _T_536 ? _GEN_235 : mem_234; // @[AsyncQueue.scala 47:24]
  assign _GEN_492 = _T_536 ? _GEN_236 : mem_235; // @[AsyncQueue.scala 47:24]
  assign _GEN_493 = _T_536 ? _GEN_237 : mem_236; // @[AsyncQueue.scala 47:24]
  assign _GEN_494 = _T_536 ? _GEN_238 : mem_237; // @[AsyncQueue.scala 47:24]
  assign _GEN_495 = _T_536 ? _GEN_239 : mem_238; // @[AsyncQueue.scala 47:24]
  assign _GEN_496 = _T_536 ? _GEN_240 : mem_239; // @[AsyncQueue.scala 47:24]
  assign _GEN_497 = _T_536 ? _GEN_241 : mem_240; // @[AsyncQueue.scala 47:24]
  assign _GEN_498 = _T_536 ? _GEN_242 : mem_241; // @[AsyncQueue.scala 47:24]
  assign _GEN_499 = _T_536 ? _GEN_243 : mem_242; // @[AsyncQueue.scala 47:24]
  assign _GEN_500 = _T_536 ? _GEN_244 : mem_243; // @[AsyncQueue.scala 47:24]
  assign _GEN_501 = _T_536 ? _GEN_245 : mem_244; // @[AsyncQueue.scala 47:24]
  assign _GEN_502 = _T_536 ? _GEN_246 : mem_245; // @[AsyncQueue.scala 47:24]
  assign _GEN_503 = _T_536 ? _GEN_247 : mem_246; // @[AsyncQueue.scala 47:24]
  assign _GEN_504 = _T_536 ? _GEN_248 : mem_247; // @[AsyncQueue.scala 47:24]
  assign _GEN_505 = _T_536 ? _GEN_249 : mem_248; // @[AsyncQueue.scala 47:24]
  assign _GEN_506 = _T_536 ? _GEN_250 : mem_249; // @[AsyncQueue.scala 47:24]
  assign _GEN_507 = _T_536 ? _GEN_251 : mem_250; // @[AsyncQueue.scala 47:24]
  assign _GEN_508 = _T_536 ? _GEN_252 : mem_251; // @[AsyncQueue.scala 47:24]
  assign _GEN_509 = _T_536 ? _GEN_253 : mem_252; // @[AsyncQueue.scala 47:24]
  assign _GEN_510 = _T_536 ? _GEN_254 : mem_253; // @[AsyncQueue.scala 47:24]
  assign _GEN_511 = _T_536 ? _GEN_255 : mem_254; // @[AsyncQueue.scala 47:24]
  assign _GEN_512 = _T_536 ? _GEN_256 : mem_255; // @[AsyncQueue.scala 47:24]
  assign ready_reg_1 = ready_reg_io_q; // @[AsyncQueue.scala 49:59]
  assign _T_558 = ready_reg_1 & sink_ready; // @[AsyncQueue.scala 50:29]
  assign _T_563 = io_sink_reset_n == 1'h0; // @[AsyncQueue.scala 62:36]
  assign _T_564 = reset | _T_563; // @[AsyncQueue.scala 62:33]
  assign io_enq_ready = _T_558;
  assign io_widx = widx_gray_io_q;
  assign io_mem_0 = mem_0;
  assign io_mem_1 = mem_1;
  assign io_mem_2 = mem_2;
  assign io_mem_3 = mem_3;
  assign io_mem_4 = mem_4;
  assign io_mem_5 = mem_5;
  assign io_mem_6 = mem_6;
  assign io_mem_7 = mem_7;
  assign io_mem_8 = mem_8;
  assign io_mem_9 = mem_9;
  assign io_mem_10 = mem_10;
  assign io_mem_11 = mem_11;
  assign io_mem_12 = mem_12;
  assign io_mem_13 = mem_13;
  assign io_mem_14 = mem_14;
  assign io_mem_15 = mem_15;
  assign io_mem_16 = mem_16;
  assign io_mem_17 = mem_17;
  assign io_mem_18 = mem_18;
  assign io_mem_19 = mem_19;
  assign io_mem_20 = mem_20;
  assign io_mem_21 = mem_21;
  assign io_mem_22 = mem_22;
  assign io_mem_23 = mem_23;
  assign io_mem_24 = mem_24;
  assign io_mem_25 = mem_25;
  assign io_mem_26 = mem_26;
  assign io_mem_27 = mem_27;
  assign io_mem_28 = mem_28;
  assign io_mem_29 = mem_29;
  assign io_mem_30 = mem_30;
  assign io_mem_31 = mem_31;
  assign io_mem_32 = mem_32;
  assign io_mem_33 = mem_33;
  assign io_mem_34 = mem_34;
  assign io_mem_35 = mem_35;
  assign io_mem_36 = mem_36;
  assign io_mem_37 = mem_37;
  assign io_mem_38 = mem_38;
  assign io_mem_39 = mem_39;
  assign io_mem_40 = mem_40;
  assign io_mem_41 = mem_41;
  assign io_mem_42 = mem_42;
  assign io_mem_43 = mem_43;
  assign io_mem_44 = mem_44;
  assign io_mem_45 = mem_45;
  assign io_mem_46 = mem_46;
  assign io_mem_47 = mem_47;
  assign io_mem_48 = mem_48;
  assign io_mem_49 = mem_49;
  assign io_mem_50 = mem_50;
  assign io_mem_51 = mem_51;
  assign io_mem_52 = mem_52;
  assign io_mem_53 = mem_53;
  assign io_mem_54 = mem_54;
  assign io_mem_55 = mem_55;
  assign io_mem_56 = mem_56;
  assign io_mem_57 = mem_57;
  assign io_mem_58 = mem_58;
  assign io_mem_59 = mem_59;
  assign io_mem_60 = mem_60;
  assign io_mem_61 = mem_61;
  assign io_mem_62 = mem_62;
  assign io_mem_63 = mem_63;
  assign io_mem_64 = mem_64;
  assign io_mem_65 = mem_65;
  assign io_mem_66 = mem_66;
  assign io_mem_67 = mem_67;
  assign io_mem_68 = mem_68;
  assign io_mem_69 = mem_69;
  assign io_mem_70 = mem_70;
  assign io_mem_71 = mem_71;
  assign io_mem_72 = mem_72;
  assign io_mem_73 = mem_73;
  assign io_mem_74 = mem_74;
  assign io_mem_75 = mem_75;
  assign io_mem_76 = mem_76;
  assign io_mem_77 = mem_77;
  assign io_mem_78 = mem_78;
  assign io_mem_79 = mem_79;
  assign io_mem_80 = mem_80;
  assign io_mem_81 = mem_81;
  assign io_mem_82 = mem_82;
  assign io_mem_83 = mem_83;
  assign io_mem_84 = mem_84;
  assign io_mem_85 = mem_85;
  assign io_mem_86 = mem_86;
  assign io_mem_87 = mem_87;
  assign io_mem_88 = mem_88;
  assign io_mem_89 = mem_89;
  assign io_mem_90 = mem_90;
  assign io_mem_91 = mem_91;
  assign io_mem_92 = mem_92;
  assign io_mem_93 = mem_93;
  assign io_mem_94 = mem_94;
  assign io_mem_95 = mem_95;
  assign io_mem_96 = mem_96;
  assign io_mem_97 = mem_97;
  assign io_mem_98 = mem_98;
  assign io_mem_99 = mem_99;
  assign io_mem_100 = mem_100;
  assign io_mem_101 = mem_101;
  assign io_mem_102 = mem_102;
  assign io_mem_103 = mem_103;
  assign io_mem_104 = mem_104;
  assign io_mem_105 = mem_105;
  assign io_mem_106 = mem_106;
  assign io_mem_107 = mem_107;
  assign io_mem_108 = mem_108;
  assign io_mem_109 = mem_109;
  assign io_mem_110 = mem_110;
  assign io_mem_111 = mem_111;
  assign io_mem_112 = mem_112;
  assign io_mem_113 = mem_113;
  assign io_mem_114 = mem_114;
  assign io_mem_115 = mem_115;
  assign io_mem_116 = mem_116;
  assign io_mem_117 = mem_117;
  assign io_mem_118 = mem_118;
  assign io_mem_119 = mem_119;
  assign io_mem_120 = mem_120;
  assign io_mem_121 = mem_121;
  assign io_mem_122 = mem_122;
  assign io_mem_123 = mem_123;
  assign io_mem_124 = mem_124;
  assign io_mem_125 = mem_125;
  assign io_mem_126 = mem_126;
  assign io_mem_127 = mem_127;
  assign io_mem_128 = mem_128;
  assign io_mem_129 = mem_129;
  assign io_mem_130 = mem_130;
  assign io_mem_131 = mem_131;
  assign io_mem_132 = mem_132;
  assign io_mem_133 = mem_133;
  assign io_mem_134 = mem_134;
  assign io_mem_135 = mem_135;
  assign io_mem_136 = mem_136;
  assign io_mem_137 = mem_137;
  assign io_mem_138 = mem_138;
  assign io_mem_139 = mem_139;
  assign io_mem_140 = mem_140;
  assign io_mem_141 = mem_141;
  assign io_mem_142 = mem_142;
  assign io_mem_143 = mem_143;
  assign io_mem_144 = mem_144;
  assign io_mem_145 = mem_145;
  assign io_mem_146 = mem_146;
  assign io_mem_147 = mem_147;
  assign io_mem_148 = mem_148;
  assign io_mem_149 = mem_149;
  assign io_mem_150 = mem_150;
  assign io_mem_151 = mem_151;
  assign io_mem_152 = mem_152;
  assign io_mem_153 = mem_153;
  assign io_mem_154 = mem_154;
  assign io_mem_155 = mem_155;
  assign io_mem_156 = mem_156;
  assign io_mem_157 = mem_157;
  assign io_mem_158 = mem_158;
  assign io_mem_159 = mem_159;
  assign io_mem_160 = mem_160;
  assign io_mem_161 = mem_161;
  assign io_mem_162 = mem_162;
  assign io_mem_163 = mem_163;
  assign io_mem_164 = mem_164;
  assign io_mem_165 = mem_165;
  assign io_mem_166 = mem_166;
  assign io_mem_167 = mem_167;
  assign io_mem_168 = mem_168;
  assign io_mem_169 = mem_169;
  assign io_mem_170 = mem_170;
  assign io_mem_171 = mem_171;
  assign io_mem_172 = mem_172;
  assign io_mem_173 = mem_173;
  assign io_mem_174 = mem_174;
  assign io_mem_175 = mem_175;
  assign io_mem_176 = mem_176;
  assign io_mem_177 = mem_177;
  assign io_mem_178 = mem_178;
  assign io_mem_179 = mem_179;
  assign io_mem_180 = mem_180;
  assign io_mem_181 = mem_181;
  assign io_mem_182 = mem_182;
  assign io_mem_183 = mem_183;
  assign io_mem_184 = mem_184;
  assign io_mem_185 = mem_185;
  assign io_mem_186 = mem_186;
  assign io_mem_187 = mem_187;
  assign io_mem_188 = mem_188;
  assign io_mem_189 = mem_189;
  assign io_mem_190 = mem_190;
  assign io_mem_191 = mem_191;
  assign io_mem_192 = mem_192;
  assign io_mem_193 = mem_193;
  assign io_mem_194 = mem_194;
  assign io_mem_195 = mem_195;
  assign io_mem_196 = mem_196;
  assign io_mem_197 = mem_197;
  assign io_mem_198 = mem_198;
  assign io_mem_199 = mem_199;
  assign io_mem_200 = mem_200;
  assign io_mem_201 = mem_201;
  assign io_mem_202 = mem_202;
  assign io_mem_203 = mem_203;
  assign io_mem_204 = mem_204;
  assign io_mem_205 = mem_205;
  assign io_mem_206 = mem_206;
  assign io_mem_207 = mem_207;
  assign io_mem_208 = mem_208;
  assign io_mem_209 = mem_209;
  assign io_mem_210 = mem_210;
  assign io_mem_211 = mem_211;
  assign io_mem_212 = mem_212;
  assign io_mem_213 = mem_213;
  assign io_mem_214 = mem_214;
  assign io_mem_215 = mem_215;
  assign io_mem_216 = mem_216;
  assign io_mem_217 = mem_217;
  assign io_mem_218 = mem_218;
  assign io_mem_219 = mem_219;
  assign io_mem_220 = mem_220;
  assign io_mem_221 = mem_221;
  assign io_mem_222 = mem_222;
  assign io_mem_223 = mem_223;
  assign io_mem_224 = mem_224;
  assign io_mem_225 = mem_225;
  assign io_mem_226 = mem_226;
  assign io_mem_227 = mem_227;
  assign io_mem_228 = mem_228;
  assign io_mem_229 = mem_229;
  assign io_mem_230 = mem_230;
  assign io_mem_231 = mem_231;
  assign io_mem_232 = mem_232;
  assign io_mem_233 = mem_233;
  assign io_mem_234 = mem_234;
  assign io_mem_235 = mem_235;
  assign io_mem_236 = mem_236;
  assign io_mem_237 = mem_237;
  assign io_mem_238 = mem_238;
  assign io_mem_239 = mem_239;
  assign io_mem_240 = mem_240;
  assign io_mem_241 = mem_241;
  assign io_mem_242 = mem_242;
  assign io_mem_243 = mem_243;
  assign io_mem_244 = mem_244;
  assign io_mem_245 = mem_245;
  assign io_mem_246 = mem_246;
  assign io_mem_247 = mem_247;
  assign io_mem_248 = mem_248;
  assign io_mem_249 = mem_249;
  assign io_mem_250 = mem_250;
  assign io_mem_251 = mem_251;
  assign io_mem_252 = mem_252;
  assign io_mem_253 = mem_253;
  assign io_mem_254 = mem_254;
  assign io_mem_255 = mem_255;
  assign io_widx_valid = AsyncValidSync_io_out;
  assign widx_bin_clock = clock;
  assign widx_bin_reset = reset;
  assign widx_bin_io_d = _T_545;
  assign widx_bin_io_en = 1'h1;
  assign ridx_gray_clock = clock;
  assign ridx_gray_reset = reset;
  assign ridx_gray_io_d = io_ridx;
  assign ready_reg_clock = clock;
  assign ready_reg_reset = reset;
  assign ready_reg_io_d = ready;
  assign ready_reg_io_en = 1'h1;
  assign widx_gray_clock = clock;
  assign widx_gray_reset = reset;
  assign widx_gray_io_d = widx;
  assign widx_gray_io_en = 1'h1;
  assign AsyncValidSync_clock = clock;
  assign AsyncValidSync_reset = _T_564;
  assign AsyncValidSync_1_clock = clock;
  assign AsyncValidSync_1_reset = _T_564;
  assign AsyncValidSync_1_io_in = io_ridx_valid;
  assign AsyncValidSync_2_clock = clock;
  assign AsyncValidSync_2_reset = reset;
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  mem_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  mem_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  mem_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  mem_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  mem_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  mem_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  mem_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  mem_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  mem_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  mem_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  mem_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  mem_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  mem_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  mem_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  mem_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  mem_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  mem_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  mem_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  mem_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  mem_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  mem_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  mem_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  mem_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  mem_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  mem_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  mem_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  mem_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  mem_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  mem_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  mem_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  mem_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  mem_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  mem_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  mem_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  mem_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  mem_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  mem_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  mem_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  mem_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  mem_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  mem_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  mem_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  mem_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  mem_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  mem_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  mem_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  mem_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  mem_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  mem_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  mem_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  mem_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  mem_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  mem_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  mem_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  mem_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  mem_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  mem_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  mem_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  mem_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  mem_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  mem_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  mem_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  mem_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  mem_64 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  mem_65 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  mem_66 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  mem_67 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  mem_68 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  mem_69 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  mem_70 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  mem_71 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  mem_72 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  mem_73 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  mem_74 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  mem_75 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  mem_76 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  mem_77 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  mem_78 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  mem_79 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  mem_80 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  mem_81 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  mem_82 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  mem_83 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  mem_84 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  mem_85 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  mem_86 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  mem_87 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  mem_88 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  mem_89 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  mem_90 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  mem_91 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  mem_92 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  mem_93 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  mem_94 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  mem_95 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  mem_96 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  mem_97 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  mem_98 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  mem_99 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  mem_100 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  mem_101 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  mem_102 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  mem_103 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  mem_104 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  mem_105 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  mem_106 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  mem_107 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  mem_108 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  mem_109 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  mem_110 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  mem_111 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  mem_112 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  mem_113 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  mem_114 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  mem_115 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  mem_116 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  mem_117 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  mem_118 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  mem_119 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  mem_120 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  mem_121 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  mem_122 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  mem_123 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  mem_124 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  mem_125 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  mem_126 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  mem_127 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  mem_128 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  mem_129 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  mem_130 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  mem_131 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  mem_132 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  mem_133 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  mem_134 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  mem_135 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  mem_136 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  mem_137 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  mem_138 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  mem_139 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  mem_140 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  mem_141 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  mem_142 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  mem_143 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  mem_144 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  mem_145 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  mem_146 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  mem_147 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  mem_148 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  mem_149 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  mem_150 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  mem_151 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  mem_152 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  mem_153 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  mem_154 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  mem_155 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  mem_156 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  mem_157 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  mem_158 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  mem_159 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  mem_160 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  mem_161 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  mem_162 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  mem_163 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  mem_164 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  mem_165 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  mem_166 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  mem_167 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  mem_168 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  mem_169 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  mem_170 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  mem_171 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  mem_172 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  mem_173 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  mem_174 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  mem_175 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  mem_176 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  mem_177 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  mem_178 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  mem_179 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  mem_180 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  mem_181 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  mem_182 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  mem_183 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  mem_184 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  mem_185 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  mem_186 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  mem_187 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  mem_188 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  mem_189 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  mem_190 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  mem_191 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  mem_192 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  mem_193 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{$random}};
  mem_194 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{$random}};
  mem_195 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{$random}};
  mem_196 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{$random}};
  mem_197 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{$random}};
  mem_198 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{$random}};
  mem_199 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{$random}};
  mem_200 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{$random}};
  mem_201 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{$random}};
  mem_202 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{$random}};
  mem_203 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{$random}};
  mem_204 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{$random}};
  mem_205 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{$random}};
  mem_206 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{$random}};
  mem_207 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{$random}};
  mem_208 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{$random}};
  mem_209 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{$random}};
  mem_210 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{$random}};
  mem_211 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{$random}};
  mem_212 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{$random}};
  mem_213 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{$random}};
  mem_214 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{$random}};
  mem_215 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{$random}};
  mem_216 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{$random}};
  mem_217 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{$random}};
  mem_218 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{$random}};
  mem_219 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{$random}};
  mem_220 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{$random}};
  mem_221 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{$random}};
  mem_222 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{$random}};
  mem_223 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{$random}};
  mem_224 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{$random}};
  mem_225 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{$random}};
  mem_226 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{$random}};
  mem_227 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{$random}};
  mem_228 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{$random}};
  mem_229 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{$random}};
  mem_230 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{$random}};
  mem_231 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{$random}};
  mem_232 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{$random}};
  mem_233 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{$random}};
  mem_234 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{$random}};
  mem_235 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{$random}};
  mem_236 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{$random}};
  mem_237 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{$random}};
  mem_238 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{$random}};
  mem_239 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{$random}};
  mem_240 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{$random}};
  mem_241 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{$random}};
  mem_242 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{$random}};
  mem_243 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{$random}};
  mem_244 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{$random}};
  mem_245 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{$random}};
  mem_246 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{$random}};
  mem_247 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{$random}};
  mem_248 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{$random}};
  mem_249 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{$random}};
  mem_250 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{$random}};
  mem_251 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{$random}};
  mem_252 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{$random}};
  mem_253 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{$random}};
  mem_254 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{$random}};
  mem_255 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_536) begin
      if (8'h0 == index) begin
        mem_0 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1 == index) begin
        mem_1 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2 == index) begin
        mem_2 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3 == index) begin
        mem_3 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4 == index) begin
        mem_4 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5 == index) begin
        mem_5 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6 == index) begin
        mem_6 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7 == index) begin
        mem_7 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8 == index) begin
        mem_8 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9 == index) begin
        mem_9 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha == index) begin
        mem_10 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb == index) begin
        mem_11 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc == index) begin
        mem_12 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd == index) begin
        mem_13 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he == index) begin
        mem_14 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf == index) begin
        mem_15 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h10 == index) begin
        mem_16 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h11 == index) begin
        mem_17 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h12 == index) begin
        mem_18 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h13 == index) begin
        mem_19 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h14 == index) begin
        mem_20 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h15 == index) begin
        mem_21 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h16 == index) begin
        mem_22 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h17 == index) begin
        mem_23 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h18 == index) begin
        mem_24 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h19 == index) begin
        mem_25 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1a == index) begin
        mem_26 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1b == index) begin
        mem_27 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1c == index) begin
        mem_28 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1d == index) begin
        mem_29 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1e == index) begin
        mem_30 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1f == index) begin
        mem_31 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h20 == index) begin
        mem_32 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h21 == index) begin
        mem_33 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h22 == index) begin
        mem_34 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h23 == index) begin
        mem_35 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h24 == index) begin
        mem_36 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h25 == index) begin
        mem_37 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h26 == index) begin
        mem_38 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h27 == index) begin
        mem_39 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h28 == index) begin
        mem_40 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h29 == index) begin
        mem_41 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2a == index) begin
        mem_42 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2b == index) begin
        mem_43 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2c == index) begin
        mem_44 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2d == index) begin
        mem_45 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2e == index) begin
        mem_46 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2f == index) begin
        mem_47 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h30 == index) begin
        mem_48 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h31 == index) begin
        mem_49 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h32 == index) begin
        mem_50 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h33 == index) begin
        mem_51 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h34 == index) begin
        mem_52 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h35 == index) begin
        mem_53 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h36 == index) begin
        mem_54 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h37 == index) begin
        mem_55 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h38 == index) begin
        mem_56 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h39 == index) begin
        mem_57 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3a == index) begin
        mem_58 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3b == index) begin
        mem_59 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3c == index) begin
        mem_60 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3d == index) begin
        mem_61 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3e == index) begin
        mem_62 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3f == index) begin
        mem_63 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h40 == index) begin
        mem_64 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h41 == index) begin
        mem_65 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h42 == index) begin
        mem_66 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h43 == index) begin
        mem_67 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h44 == index) begin
        mem_68 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h45 == index) begin
        mem_69 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h46 == index) begin
        mem_70 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h47 == index) begin
        mem_71 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h48 == index) begin
        mem_72 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h49 == index) begin
        mem_73 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4a == index) begin
        mem_74 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4b == index) begin
        mem_75 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4c == index) begin
        mem_76 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4d == index) begin
        mem_77 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4e == index) begin
        mem_78 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4f == index) begin
        mem_79 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h50 == index) begin
        mem_80 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h51 == index) begin
        mem_81 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h52 == index) begin
        mem_82 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h53 == index) begin
        mem_83 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h54 == index) begin
        mem_84 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h55 == index) begin
        mem_85 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h56 == index) begin
        mem_86 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h57 == index) begin
        mem_87 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h58 == index) begin
        mem_88 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h59 == index) begin
        mem_89 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5a == index) begin
        mem_90 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5b == index) begin
        mem_91 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5c == index) begin
        mem_92 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5d == index) begin
        mem_93 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5e == index) begin
        mem_94 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5f == index) begin
        mem_95 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h60 == index) begin
        mem_96 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h61 == index) begin
        mem_97 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h62 == index) begin
        mem_98 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h63 == index) begin
        mem_99 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h64 == index) begin
        mem_100 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h65 == index) begin
        mem_101 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h66 == index) begin
        mem_102 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h67 == index) begin
        mem_103 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h68 == index) begin
        mem_104 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h69 == index) begin
        mem_105 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6a == index) begin
        mem_106 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6b == index) begin
        mem_107 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6c == index) begin
        mem_108 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6d == index) begin
        mem_109 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6e == index) begin
        mem_110 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6f == index) begin
        mem_111 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h70 == index) begin
        mem_112 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h71 == index) begin
        mem_113 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h72 == index) begin
        mem_114 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h73 == index) begin
        mem_115 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h74 == index) begin
        mem_116 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h75 == index) begin
        mem_117 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h76 == index) begin
        mem_118 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h77 == index) begin
        mem_119 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h78 == index) begin
        mem_120 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h79 == index) begin
        mem_121 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7a == index) begin
        mem_122 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7b == index) begin
        mem_123 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7c == index) begin
        mem_124 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7d == index) begin
        mem_125 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7e == index) begin
        mem_126 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7f == index) begin
        mem_127 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h80 == index) begin
        mem_128 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h81 == index) begin
        mem_129 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h82 == index) begin
        mem_130 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h83 == index) begin
        mem_131 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h84 == index) begin
        mem_132 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h85 == index) begin
        mem_133 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h86 == index) begin
        mem_134 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h87 == index) begin
        mem_135 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h88 == index) begin
        mem_136 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h89 == index) begin
        mem_137 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8a == index) begin
        mem_138 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8b == index) begin
        mem_139 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8c == index) begin
        mem_140 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8d == index) begin
        mem_141 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8e == index) begin
        mem_142 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8f == index) begin
        mem_143 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h90 == index) begin
        mem_144 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h91 == index) begin
        mem_145 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h92 == index) begin
        mem_146 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h93 == index) begin
        mem_147 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h94 == index) begin
        mem_148 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h95 == index) begin
        mem_149 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h96 == index) begin
        mem_150 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h97 == index) begin
        mem_151 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h98 == index) begin
        mem_152 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h99 == index) begin
        mem_153 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9a == index) begin
        mem_154 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9b == index) begin
        mem_155 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9c == index) begin
        mem_156 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9d == index) begin
        mem_157 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9e == index) begin
        mem_158 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9f == index) begin
        mem_159 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha0 == index) begin
        mem_160 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha1 == index) begin
        mem_161 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha2 == index) begin
        mem_162 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha3 == index) begin
        mem_163 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha4 == index) begin
        mem_164 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha5 == index) begin
        mem_165 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha6 == index) begin
        mem_166 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha7 == index) begin
        mem_167 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha8 == index) begin
        mem_168 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha9 == index) begin
        mem_169 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'haa == index) begin
        mem_170 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hab == index) begin
        mem_171 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hac == index) begin
        mem_172 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'had == index) begin
        mem_173 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hae == index) begin
        mem_174 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'haf == index) begin
        mem_175 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb0 == index) begin
        mem_176 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb1 == index) begin
        mem_177 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb2 == index) begin
        mem_178 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb3 == index) begin
        mem_179 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb4 == index) begin
        mem_180 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb5 == index) begin
        mem_181 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb6 == index) begin
        mem_182 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb7 == index) begin
        mem_183 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb8 == index) begin
        mem_184 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb9 == index) begin
        mem_185 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hba == index) begin
        mem_186 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hbb == index) begin
        mem_187 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hbc == index) begin
        mem_188 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hbd == index) begin
        mem_189 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hbe == index) begin
        mem_190 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hbf == index) begin
        mem_191 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc0 == index) begin
        mem_192 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc1 == index) begin
        mem_193 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc2 == index) begin
        mem_194 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc3 == index) begin
        mem_195 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc4 == index) begin
        mem_196 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc5 == index) begin
        mem_197 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc6 == index) begin
        mem_198 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc7 == index) begin
        mem_199 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc8 == index) begin
        mem_200 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc9 == index) begin
        mem_201 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hca == index) begin
        mem_202 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hcb == index) begin
        mem_203 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hcc == index) begin
        mem_204 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hcd == index) begin
        mem_205 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hce == index) begin
        mem_206 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hcf == index) begin
        mem_207 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd0 == index) begin
        mem_208 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd1 == index) begin
        mem_209 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd2 == index) begin
        mem_210 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd3 == index) begin
        mem_211 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd4 == index) begin
        mem_212 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd5 == index) begin
        mem_213 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd6 == index) begin
        mem_214 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd7 == index) begin
        mem_215 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd8 == index) begin
        mem_216 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd9 == index) begin
        mem_217 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hda == index) begin
        mem_218 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hdb == index) begin
        mem_219 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hdc == index) begin
        mem_220 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hdd == index) begin
        mem_221 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hde == index) begin
        mem_222 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hdf == index) begin
        mem_223 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he0 == index) begin
        mem_224 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he1 == index) begin
        mem_225 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he2 == index) begin
        mem_226 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he3 == index) begin
        mem_227 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he4 == index) begin
        mem_228 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he5 == index) begin
        mem_229 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he6 == index) begin
        mem_230 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he7 == index) begin
        mem_231 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he8 == index) begin
        mem_232 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he9 == index) begin
        mem_233 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hea == index) begin
        mem_234 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'heb == index) begin
        mem_235 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hec == index) begin
        mem_236 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hed == index) begin
        mem_237 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hee == index) begin
        mem_238 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hef == index) begin
        mem_239 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf0 == index) begin
        mem_240 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf1 == index) begin
        mem_241 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf2 == index) begin
        mem_242 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf3 == index) begin
        mem_243 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf4 == index) begin
        mem_244 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf5 == index) begin
        mem_245 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf6 == index) begin
        mem_246 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf7 == index) begin
        mem_247 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf8 == index) begin
        mem_248 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf9 == index) begin
        mem_249 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hfa == index) begin
        mem_250 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hfb == index) begin
        mem_251 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hfc == index) begin
        mem_252 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hfd == index) begin
        mem_253 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hfe == index) begin
        mem_254 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hff == index) begin
        mem_255 <= io_enq_bits;
      end
    end
  end
endmodule
module SynchronizerShiftReg_w1_d1(
  input   clock,
  input   io_d,
  output  io_q
);
  reg  sync_0; // @[ShiftReg.scala 114:16]
  reg [31:0] _RAND_0;
  assign io_q = sync_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  sync_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    sync_0 <= io_d;
  end
endmodule
module AsyncValidSync_3(
  input   clock,
  input   reset,
  output  io_out
);
  wire  sink_valid_clock; // @[ShiftReg.scala 47:23]
  wire  sink_valid_reset; // @[ShiftReg.scala 47:23]
  wire  sink_valid_io_q; // @[ShiftReg.scala 47:23]
  wire  _T_5; // @[ShiftReg.scala 50:24]
  AsyncResetSynchronizerShiftReg_w1_d4_i0 sink_valid ( // @[ShiftReg.scala 47:23]
    .clock(sink_valid_clock),
    .reset(sink_valid_reset),
    .io_q(sink_valid_io_q)
  );
  assign _T_5 = sink_valid_io_q; // @[ShiftReg.scala 50:24]
  assign io_out = _T_5;
  assign sink_valid_clock = clock;
  assign sink_valid_reset = reset;
endmodule
module AsyncValidSync_4(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  source_extend_clock; // @[ShiftReg.scala 47:23]
  wire  source_extend_reset; // @[ShiftReg.scala 47:23]
  wire  source_extend_io_d; // @[ShiftReg.scala 47:23]
  wire  source_extend_io_q; // @[ShiftReg.scala 47:23]
  wire  _T_5; // @[ShiftReg.scala 50:24]
  AsyncResetSynchronizerShiftReg_w1_d1_i0 source_extend ( // @[ShiftReg.scala 47:23]
    .clock(source_extend_clock),
    .reset(source_extend_reset),
    .io_d(source_extend_io_d),
    .io_q(source_extend_io_q)
  );
  assign _T_5 = source_extend_io_q; // @[ShiftReg.scala 50:24]
  assign io_out = _T_5;
  assign source_extend_clock = clock;
  assign source_extend_reset = reset;
  assign source_extend_io_d = io_in;
endmodule
module AsyncValidSync_5(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  source_valid_clock; // @[ShiftReg.scala 47:23]
  wire  source_valid_reset; // @[ShiftReg.scala 47:23]
  wire  source_valid_io_d; // @[ShiftReg.scala 47:23]
  wire  source_valid_io_q; // @[ShiftReg.scala 47:23]
  wire  _T_5; // @[ShiftReg.scala 50:24]
  AsyncResetSynchronizerShiftReg_w1_d3_i0 source_valid ( // @[ShiftReg.scala 47:23]
    .clock(source_valid_clock),
    .reset(source_valid_reset),
    .io_d(source_valid_io_d),
    .io_q(source_valid_io_q)
  );
  assign _T_5 = source_valid_io_q; // @[ShiftReg.scala 50:24]
  assign io_out = _T_5;
  assign source_valid_clock = clock;
  assign source_valid_reset = reset;
  assign source_valid_io_d = io_in;
endmodule
module AsyncQueueSink(
  input        clock,
  input        reset,
  input        io_deq_ready,
  output       io_deq_valid,
  output       io_deq_bits,
  output [8:0] io_ridx,
  input  [8:0] io_widx,
  input        io_mem_0,
  input        io_mem_1,
  input        io_mem_2,
  input        io_mem_3,
  input        io_mem_4,
  input        io_mem_5,
  input        io_mem_6,
  input        io_mem_7,
  input        io_mem_8,
  input        io_mem_9,
  input        io_mem_10,
  input        io_mem_11,
  input        io_mem_12,
  input        io_mem_13,
  input        io_mem_14,
  input        io_mem_15,
  input        io_mem_16,
  input        io_mem_17,
  input        io_mem_18,
  input        io_mem_19,
  input        io_mem_20,
  input        io_mem_21,
  input        io_mem_22,
  input        io_mem_23,
  input        io_mem_24,
  input        io_mem_25,
  input        io_mem_26,
  input        io_mem_27,
  input        io_mem_28,
  input        io_mem_29,
  input        io_mem_30,
  input        io_mem_31,
  input        io_mem_32,
  input        io_mem_33,
  input        io_mem_34,
  input        io_mem_35,
  input        io_mem_36,
  input        io_mem_37,
  input        io_mem_38,
  input        io_mem_39,
  input        io_mem_40,
  input        io_mem_41,
  input        io_mem_42,
  input        io_mem_43,
  input        io_mem_44,
  input        io_mem_45,
  input        io_mem_46,
  input        io_mem_47,
  input        io_mem_48,
  input        io_mem_49,
  input        io_mem_50,
  input        io_mem_51,
  input        io_mem_52,
  input        io_mem_53,
  input        io_mem_54,
  input        io_mem_55,
  input        io_mem_56,
  input        io_mem_57,
  input        io_mem_58,
  input        io_mem_59,
  input        io_mem_60,
  input        io_mem_61,
  input        io_mem_62,
  input        io_mem_63,
  input        io_mem_64,
  input        io_mem_65,
  input        io_mem_66,
  input        io_mem_67,
  input        io_mem_68,
  input        io_mem_69,
  input        io_mem_70,
  input        io_mem_71,
  input        io_mem_72,
  input        io_mem_73,
  input        io_mem_74,
  input        io_mem_75,
  input        io_mem_76,
  input        io_mem_77,
  input        io_mem_78,
  input        io_mem_79,
  input        io_mem_80,
  input        io_mem_81,
  input        io_mem_82,
  input        io_mem_83,
  input        io_mem_84,
  input        io_mem_85,
  input        io_mem_86,
  input        io_mem_87,
  input        io_mem_88,
  input        io_mem_89,
  input        io_mem_90,
  input        io_mem_91,
  input        io_mem_92,
  input        io_mem_93,
  input        io_mem_94,
  input        io_mem_95,
  input        io_mem_96,
  input        io_mem_97,
  input        io_mem_98,
  input        io_mem_99,
  input        io_mem_100,
  input        io_mem_101,
  input        io_mem_102,
  input        io_mem_103,
  input        io_mem_104,
  input        io_mem_105,
  input        io_mem_106,
  input        io_mem_107,
  input        io_mem_108,
  input        io_mem_109,
  input        io_mem_110,
  input        io_mem_111,
  input        io_mem_112,
  input        io_mem_113,
  input        io_mem_114,
  input        io_mem_115,
  input        io_mem_116,
  input        io_mem_117,
  input        io_mem_118,
  input        io_mem_119,
  input        io_mem_120,
  input        io_mem_121,
  input        io_mem_122,
  input        io_mem_123,
  input        io_mem_124,
  input        io_mem_125,
  input        io_mem_126,
  input        io_mem_127,
  input        io_mem_128,
  input        io_mem_129,
  input        io_mem_130,
  input        io_mem_131,
  input        io_mem_132,
  input        io_mem_133,
  input        io_mem_134,
  input        io_mem_135,
  input        io_mem_136,
  input        io_mem_137,
  input        io_mem_138,
  input        io_mem_139,
  input        io_mem_140,
  input        io_mem_141,
  input        io_mem_142,
  input        io_mem_143,
  input        io_mem_144,
  input        io_mem_145,
  input        io_mem_146,
  input        io_mem_147,
  input        io_mem_148,
  input        io_mem_149,
  input        io_mem_150,
  input        io_mem_151,
  input        io_mem_152,
  input        io_mem_153,
  input        io_mem_154,
  input        io_mem_155,
  input        io_mem_156,
  input        io_mem_157,
  input        io_mem_158,
  input        io_mem_159,
  input        io_mem_160,
  input        io_mem_161,
  input        io_mem_162,
  input        io_mem_163,
  input        io_mem_164,
  input        io_mem_165,
  input        io_mem_166,
  input        io_mem_167,
  input        io_mem_168,
  input        io_mem_169,
  input        io_mem_170,
  input        io_mem_171,
  input        io_mem_172,
  input        io_mem_173,
  input        io_mem_174,
  input        io_mem_175,
  input        io_mem_176,
  input        io_mem_177,
  input        io_mem_178,
  input        io_mem_179,
  input        io_mem_180,
  input        io_mem_181,
  input        io_mem_182,
  input        io_mem_183,
  input        io_mem_184,
  input        io_mem_185,
  input        io_mem_186,
  input        io_mem_187,
  input        io_mem_188,
  input        io_mem_189,
  input        io_mem_190,
  input        io_mem_191,
  input        io_mem_192,
  input        io_mem_193,
  input        io_mem_194,
  input        io_mem_195,
  input        io_mem_196,
  input        io_mem_197,
  input        io_mem_198,
  input        io_mem_199,
  input        io_mem_200,
  input        io_mem_201,
  input        io_mem_202,
  input        io_mem_203,
  input        io_mem_204,
  input        io_mem_205,
  input        io_mem_206,
  input        io_mem_207,
  input        io_mem_208,
  input        io_mem_209,
  input        io_mem_210,
  input        io_mem_211,
  input        io_mem_212,
  input        io_mem_213,
  input        io_mem_214,
  input        io_mem_215,
  input        io_mem_216,
  input        io_mem_217,
  input        io_mem_218,
  input        io_mem_219,
  input        io_mem_220,
  input        io_mem_221,
  input        io_mem_222,
  input        io_mem_223,
  input        io_mem_224,
  input        io_mem_225,
  input        io_mem_226,
  input        io_mem_227,
  input        io_mem_228,
  input        io_mem_229,
  input        io_mem_230,
  input        io_mem_231,
  input        io_mem_232,
  input        io_mem_233,
  input        io_mem_234,
  input        io_mem_235,
  input        io_mem_236,
  input        io_mem_237,
  input        io_mem_238,
  input        io_mem_239,
  input        io_mem_240,
  input        io_mem_241,
  input        io_mem_242,
  input        io_mem_243,
  input        io_mem_244,
  input        io_mem_245,
  input        io_mem_246,
  input        io_mem_247,
  input        io_mem_248,
  input        io_mem_249,
  input        io_mem_250,
  input        io_mem_251,
  input        io_mem_252,
  input        io_mem_253,
  input        io_mem_254,
  input        io_mem_255,
  input        io_source_reset_n,
  output       io_ridx_valid,
  input        io_widx_valid
);
  wire  ridx_bin_clock; // @[AsyncResetReg.scala 110:21]
  wire  ridx_bin_reset; // @[AsyncResetReg.scala 110:21]
  wire [8:0] ridx_bin_io_d; // @[AsyncResetReg.scala 110:21]
  wire [8:0] ridx_bin_io_q; // @[AsyncResetReg.scala 110:21]
  wire  ridx_bin_io_en; // @[AsyncResetReg.scala 110:21]
  wire  widx_gray_clock; // @[ShiftReg.scala 47:23]
  wire  widx_gray_reset; // @[ShiftReg.scala 47:23]
  wire [8:0] widx_gray_io_d; // @[ShiftReg.scala 47:23]
  wire [8:0] widx_gray_io_q; // @[ShiftReg.scala 47:23]
  wire  deq_bits_reg_clock; // @[ShiftReg.scala 47:23]
  wire  deq_bits_reg_io_d; // @[ShiftReg.scala 47:23]
  wire  deq_bits_reg_io_q; // @[ShiftReg.scala 47:23]
  wire  valid_reg_clock; // @[AsyncResetReg.scala 110:21]
  wire  valid_reg_reset; // @[AsyncResetReg.scala 110:21]
  wire  valid_reg_io_d; // @[AsyncResetReg.scala 110:21]
  wire  valid_reg_io_q; // @[AsyncResetReg.scala 110:21]
  wire  valid_reg_io_en; // @[AsyncResetReg.scala 110:21]
  wire  ridx_gray_clock; // @[AsyncResetReg.scala 110:21]
  wire  ridx_gray_reset; // @[AsyncResetReg.scala 110:21]
  wire [8:0] ridx_gray_io_d; // @[AsyncResetReg.scala 110:21]
  wire [8:0] ridx_gray_io_q; // @[AsyncResetReg.scala 110:21]
  wire  ridx_gray_io_en; // @[AsyncResetReg.scala 110:21]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 124:31]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 124:31]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 124:31]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 125:31]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 125:31]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 125:31]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 125:31]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 126:31]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 126:31]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 126:31]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 126:31]
  wire  AsyncResetRegVec_w1_i0_clock; // @[AsyncResetReg.scala 110:21]
  wire  AsyncResetRegVec_w1_i0_reset; // @[AsyncResetReg.scala 110:21]
  wire  AsyncResetRegVec_w1_i0_io_d; // @[AsyncResetReg.scala 110:21]
  wire  AsyncResetRegVec_w1_i0_io_q; // @[AsyncResetReg.scala 110:21]
  wire  AsyncResetRegVec_w1_i0_io_en; // @[AsyncResetReg.scala 110:21]
  wire  _T_272; // @[Decoupled.scala 30:37]
  wire  source_ready;
  wire  _T_274; // @[AsyncQueue.scala 99:49]
  wire [8:0] _GEN_256; // @[AsyncQueue.scala 11:47]
  wire [9:0] _T_279; // @[AsyncQueue.scala 11:47]
  wire [8:0] _T_280; // @[AsyncQueue.scala 11:47]
  wire [8:0] _T_281; // @[AsyncQueue.scala 11:23]
  wire [8:0] _T_283; // @[AsyncQueue.scala 12:32]
  wire [8:0] ridx; // @[AsyncQueue.scala 12:17]
  wire [8:0] widx; // @[ShiftReg.scala 50:24]
  wire  _T_285; // @[AsyncQueue.scala 101:36]
  wire  valid; // @[AsyncQueue.scala 101:28]
  wire [7:0] _T_286; // @[AsyncQueue.scala 107:48]
  wire  _T_287; // @[AsyncQueue.scala 107:67]
  wire [7:0] _GEN_257; // @[AsyncQueue.scala 107:80]
  wire [7:0] _T_288; // @[AsyncQueue.scala 107:80]
  wire [7:0] index; // @[AsyncQueue.scala 107:60]
  wire  _GEN_1; // @[AsyncQueue.scala 113:25]
  wire  _GEN_2; // @[AsyncQueue.scala 113:25]
  wire  _GEN_3; // @[AsyncQueue.scala 113:25]
  wire  _GEN_4; // @[AsyncQueue.scala 113:25]
  wire  _GEN_5; // @[AsyncQueue.scala 113:25]
  wire  _GEN_6; // @[AsyncQueue.scala 113:25]
  wire  _GEN_7; // @[AsyncQueue.scala 113:25]
  wire  _GEN_8; // @[AsyncQueue.scala 113:25]
  wire  _GEN_9; // @[AsyncQueue.scala 113:25]
  wire  _GEN_10; // @[AsyncQueue.scala 113:25]
  wire  _GEN_11; // @[AsyncQueue.scala 113:25]
  wire  _GEN_12; // @[AsyncQueue.scala 113:25]
  wire  _GEN_13; // @[AsyncQueue.scala 113:25]
  wire  _GEN_14; // @[AsyncQueue.scala 113:25]
  wire  _GEN_15; // @[AsyncQueue.scala 113:25]
  wire  _GEN_16; // @[AsyncQueue.scala 113:25]
  wire  _GEN_17; // @[AsyncQueue.scala 113:25]
  wire  _GEN_18; // @[AsyncQueue.scala 113:25]
  wire  _GEN_19; // @[AsyncQueue.scala 113:25]
  wire  _GEN_20; // @[AsyncQueue.scala 113:25]
  wire  _GEN_21; // @[AsyncQueue.scala 113:25]
  wire  _GEN_22; // @[AsyncQueue.scala 113:25]
  wire  _GEN_23; // @[AsyncQueue.scala 113:25]
  wire  _GEN_24; // @[AsyncQueue.scala 113:25]
  wire  _GEN_25; // @[AsyncQueue.scala 113:25]
  wire  _GEN_26; // @[AsyncQueue.scala 113:25]
  wire  _GEN_27; // @[AsyncQueue.scala 113:25]
  wire  _GEN_28; // @[AsyncQueue.scala 113:25]
  wire  _GEN_29; // @[AsyncQueue.scala 113:25]
  wire  _GEN_30; // @[AsyncQueue.scala 113:25]
  wire  _GEN_31; // @[AsyncQueue.scala 113:25]
  wire  _GEN_32; // @[AsyncQueue.scala 113:25]
  wire  _GEN_33; // @[AsyncQueue.scala 113:25]
  wire  _GEN_34; // @[AsyncQueue.scala 113:25]
  wire  _GEN_35; // @[AsyncQueue.scala 113:25]
  wire  _GEN_36; // @[AsyncQueue.scala 113:25]
  wire  _GEN_37; // @[AsyncQueue.scala 113:25]
  wire  _GEN_38; // @[AsyncQueue.scala 113:25]
  wire  _GEN_39; // @[AsyncQueue.scala 113:25]
  wire  _GEN_40; // @[AsyncQueue.scala 113:25]
  wire  _GEN_41; // @[AsyncQueue.scala 113:25]
  wire  _GEN_42; // @[AsyncQueue.scala 113:25]
  wire  _GEN_43; // @[AsyncQueue.scala 113:25]
  wire  _GEN_44; // @[AsyncQueue.scala 113:25]
  wire  _GEN_45; // @[AsyncQueue.scala 113:25]
  wire  _GEN_46; // @[AsyncQueue.scala 113:25]
  wire  _GEN_47; // @[AsyncQueue.scala 113:25]
  wire  _GEN_48; // @[AsyncQueue.scala 113:25]
  wire  _GEN_49; // @[AsyncQueue.scala 113:25]
  wire  _GEN_50; // @[AsyncQueue.scala 113:25]
  wire  _GEN_51; // @[AsyncQueue.scala 113:25]
  wire  _GEN_52; // @[AsyncQueue.scala 113:25]
  wire  _GEN_53; // @[AsyncQueue.scala 113:25]
  wire  _GEN_54; // @[AsyncQueue.scala 113:25]
  wire  _GEN_55; // @[AsyncQueue.scala 113:25]
  wire  _GEN_56; // @[AsyncQueue.scala 113:25]
  wire  _GEN_57; // @[AsyncQueue.scala 113:25]
  wire  _GEN_58; // @[AsyncQueue.scala 113:25]
  wire  _GEN_59; // @[AsyncQueue.scala 113:25]
  wire  _GEN_60; // @[AsyncQueue.scala 113:25]
  wire  _GEN_61; // @[AsyncQueue.scala 113:25]
  wire  _GEN_62; // @[AsyncQueue.scala 113:25]
  wire  _GEN_63; // @[AsyncQueue.scala 113:25]
  wire  _GEN_64; // @[AsyncQueue.scala 113:25]
  wire  _GEN_65; // @[AsyncQueue.scala 113:25]
  wire  _GEN_66; // @[AsyncQueue.scala 113:25]
  wire  _GEN_67; // @[AsyncQueue.scala 113:25]
  wire  _GEN_68; // @[AsyncQueue.scala 113:25]
  wire  _GEN_69; // @[AsyncQueue.scala 113:25]
  wire  _GEN_70; // @[AsyncQueue.scala 113:25]
  wire  _GEN_71; // @[AsyncQueue.scala 113:25]
  wire  _GEN_72; // @[AsyncQueue.scala 113:25]
  wire  _GEN_73; // @[AsyncQueue.scala 113:25]
  wire  _GEN_74; // @[AsyncQueue.scala 113:25]
  wire  _GEN_75; // @[AsyncQueue.scala 113:25]
  wire  _GEN_76; // @[AsyncQueue.scala 113:25]
  wire  _GEN_77; // @[AsyncQueue.scala 113:25]
  wire  _GEN_78; // @[AsyncQueue.scala 113:25]
  wire  _GEN_79; // @[AsyncQueue.scala 113:25]
  wire  _GEN_80; // @[AsyncQueue.scala 113:25]
  wire  _GEN_81; // @[AsyncQueue.scala 113:25]
  wire  _GEN_82; // @[AsyncQueue.scala 113:25]
  wire  _GEN_83; // @[AsyncQueue.scala 113:25]
  wire  _GEN_84; // @[AsyncQueue.scala 113:25]
  wire  _GEN_85; // @[AsyncQueue.scala 113:25]
  wire  _GEN_86; // @[AsyncQueue.scala 113:25]
  wire  _GEN_87; // @[AsyncQueue.scala 113:25]
  wire  _GEN_88; // @[AsyncQueue.scala 113:25]
  wire  _GEN_89; // @[AsyncQueue.scala 113:25]
  wire  _GEN_90; // @[AsyncQueue.scala 113:25]
  wire  _GEN_91; // @[AsyncQueue.scala 113:25]
  wire  _GEN_92; // @[AsyncQueue.scala 113:25]
  wire  _GEN_93; // @[AsyncQueue.scala 113:25]
  wire  _GEN_94; // @[AsyncQueue.scala 113:25]
  wire  _GEN_95; // @[AsyncQueue.scala 113:25]
  wire  _GEN_96; // @[AsyncQueue.scala 113:25]
  wire  _GEN_97; // @[AsyncQueue.scala 113:25]
  wire  _GEN_98; // @[AsyncQueue.scala 113:25]
  wire  _GEN_99; // @[AsyncQueue.scala 113:25]
  wire  _GEN_100; // @[AsyncQueue.scala 113:25]
  wire  _GEN_101; // @[AsyncQueue.scala 113:25]
  wire  _GEN_102; // @[AsyncQueue.scala 113:25]
  wire  _GEN_103; // @[AsyncQueue.scala 113:25]
  wire  _GEN_104; // @[AsyncQueue.scala 113:25]
  wire  _GEN_105; // @[AsyncQueue.scala 113:25]
  wire  _GEN_106; // @[AsyncQueue.scala 113:25]
  wire  _GEN_107; // @[AsyncQueue.scala 113:25]
  wire  _GEN_108; // @[AsyncQueue.scala 113:25]
  wire  _GEN_109; // @[AsyncQueue.scala 113:25]
  wire  _GEN_110; // @[AsyncQueue.scala 113:25]
  wire  _GEN_111; // @[AsyncQueue.scala 113:25]
  wire  _GEN_112; // @[AsyncQueue.scala 113:25]
  wire  _GEN_113; // @[AsyncQueue.scala 113:25]
  wire  _GEN_114; // @[AsyncQueue.scala 113:25]
  wire  _GEN_115; // @[AsyncQueue.scala 113:25]
  wire  _GEN_116; // @[AsyncQueue.scala 113:25]
  wire  _GEN_117; // @[AsyncQueue.scala 113:25]
  wire  _GEN_118; // @[AsyncQueue.scala 113:25]
  wire  _GEN_119; // @[AsyncQueue.scala 113:25]
  wire  _GEN_120; // @[AsyncQueue.scala 113:25]
  wire  _GEN_121; // @[AsyncQueue.scala 113:25]
  wire  _GEN_122; // @[AsyncQueue.scala 113:25]
  wire  _GEN_123; // @[AsyncQueue.scala 113:25]
  wire  _GEN_124; // @[AsyncQueue.scala 113:25]
  wire  _GEN_125; // @[AsyncQueue.scala 113:25]
  wire  _GEN_126; // @[AsyncQueue.scala 113:25]
  wire  _GEN_127; // @[AsyncQueue.scala 113:25]
  wire  _GEN_128; // @[AsyncQueue.scala 113:25]
  wire  _GEN_129; // @[AsyncQueue.scala 113:25]
  wire  _GEN_130; // @[AsyncQueue.scala 113:25]
  wire  _GEN_131; // @[AsyncQueue.scala 113:25]
  wire  _GEN_132; // @[AsyncQueue.scala 113:25]
  wire  _GEN_133; // @[AsyncQueue.scala 113:25]
  wire  _GEN_134; // @[AsyncQueue.scala 113:25]
  wire  _GEN_135; // @[AsyncQueue.scala 113:25]
  wire  _GEN_136; // @[AsyncQueue.scala 113:25]
  wire  _GEN_137; // @[AsyncQueue.scala 113:25]
  wire  _GEN_138; // @[AsyncQueue.scala 113:25]
  wire  _GEN_139; // @[AsyncQueue.scala 113:25]
  wire  _GEN_140; // @[AsyncQueue.scala 113:25]
  wire  _GEN_141; // @[AsyncQueue.scala 113:25]
  wire  _GEN_142; // @[AsyncQueue.scala 113:25]
  wire  _GEN_143; // @[AsyncQueue.scala 113:25]
  wire  _GEN_144; // @[AsyncQueue.scala 113:25]
  wire  _GEN_145; // @[AsyncQueue.scala 113:25]
  wire  _GEN_146; // @[AsyncQueue.scala 113:25]
  wire  _GEN_147; // @[AsyncQueue.scala 113:25]
  wire  _GEN_148; // @[AsyncQueue.scala 113:25]
  wire  _GEN_149; // @[AsyncQueue.scala 113:25]
  wire  _GEN_150; // @[AsyncQueue.scala 113:25]
  wire  _GEN_151; // @[AsyncQueue.scala 113:25]
  wire  _GEN_152; // @[AsyncQueue.scala 113:25]
  wire  _GEN_153; // @[AsyncQueue.scala 113:25]
  wire  _GEN_154; // @[AsyncQueue.scala 113:25]
  wire  _GEN_155; // @[AsyncQueue.scala 113:25]
  wire  _GEN_156; // @[AsyncQueue.scala 113:25]
  wire  _GEN_157; // @[AsyncQueue.scala 113:25]
  wire  _GEN_158; // @[AsyncQueue.scala 113:25]
  wire  _GEN_159; // @[AsyncQueue.scala 113:25]
  wire  _GEN_160; // @[AsyncQueue.scala 113:25]
  wire  _GEN_161; // @[AsyncQueue.scala 113:25]
  wire  _GEN_162; // @[AsyncQueue.scala 113:25]
  wire  _GEN_163; // @[AsyncQueue.scala 113:25]
  wire  _GEN_164; // @[AsyncQueue.scala 113:25]
  wire  _GEN_165; // @[AsyncQueue.scala 113:25]
  wire  _GEN_166; // @[AsyncQueue.scala 113:25]
  wire  _GEN_167; // @[AsyncQueue.scala 113:25]
  wire  _GEN_168; // @[AsyncQueue.scala 113:25]
  wire  _GEN_169; // @[AsyncQueue.scala 113:25]
  wire  _GEN_170; // @[AsyncQueue.scala 113:25]
  wire  _GEN_171; // @[AsyncQueue.scala 113:25]
  wire  _GEN_172; // @[AsyncQueue.scala 113:25]
  wire  _GEN_173; // @[AsyncQueue.scala 113:25]
  wire  _GEN_174; // @[AsyncQueue.scala 113:25]
  wire  _GEN_175; // @[AsyncQueue.scala 113:25]
  wire  _GEN_176; // @[AsyncQueue.scala 113:25]
  wire  _GEN_177; // @[AsyncQueue.scala 113:25]
  wire  _GEN_178; // @[AsyncQueue.scala 113:25]
  wire  _GEN_179; // @[AsyncQueue.scala 113:25]
  wire  _GEN_180; // @[AsyncQueue.scala 113:25]
  wire  _GEN_181; // @[AsyncQueue.scala 113:25]
  wire  _GEN_182; // @[AsyncQueue.scala 113:25]
  wire  _GEN_183; // @[AsyncQueue.scala 113:25]
  wire  _GEN_184; // @[AsyncQueue.scala 113:25]
  wire  _GEN_185; // @[AsyncQueue.scala 113:25]
  wire  _GEN_186; // @[AsyncQueue.scala 113:25]
  wire  _GEN_187; // @[AsyncQueue.scala 113:25]
  wire  _GEN_188; // @[AsyncQueue.scala 113:25]
  wire  _GEN_189; // @[AsyncQueue.scala 113:25]
  wire  _GEN_190; // @[AsyncQueue.scala 113:25]
  wire  _GEN_191; // @[AsyncQueue.scala 113:25]
  wire  _GEN_192; // @[AsyncQueue.scala 113:25]
  wire  _GEN_193; // @[AsyncQueue.scala 113:25]
  wire  _GEN_194; // @[AsyncQueue.scala 113:25]
  wire  _GEN_195; // @[AsyncQueue.scala 113:25]
  wire  _GEN_196; // @[AsyncQueue.scala 113:25]
  wire  _GEN_197; // @[AsyncQueue.scala 113:25]
  wire  _GEN_198; // @[AsyncQueue.scala 113:25]
  wire  _GEN_199; // @[AsyncQueue.scala 113:25]
  wire  _GEN_200; // @[AsyncQueue.scala 113:25]
  wire  _GEN_201; // @[AsyncQueue.scala 113:25]
  wire  _GEN_202; // @[AsyncQueue.scala 113:25]
  wire  _GEN_203; // @[AsyncQueue.scala 113:25]
  wire  _GEN_204; // @[AsyncQueue.scala 113:25]
  wire  _GEN_205; // @[AsyncQueue.scala 113:25]
  wire  _GEN_206; // @[AsyncQueue.scala 113:25]
  wire  _GEN_207; // @[AsyncQueue.scala 113:25]
  wire  _GEN_208; // @[AsyncQueue.scala 113:25]
  wire  _GEN_209; // @[AsyncQueue.scala 113:25]
  wire  _GEN_210; // @[AsyncQueue.scala 113:25]
  wire  _GEN_211; // @[AsyncQueue.scala 113:25]
  wire  _GEN_212; // @[AsyncQueue.scala 113:25]
  wire  _GEN_213; // @[AsyncQueue.scala 113:25]
  wire  _GEN_214; // @[AsyncQueue.scala 113:25]
  wire  _GEN_215; // @[AsyncQueue.scala 113:25]
  wire  _GEN_216; // @[AsyncQueue.scala 113:25]
  wire  _GEN_217; // @[AsyncQueue.scala 113:25]
  wire  _GEN_218; // @[AsyncQueue.scala 113:25]
  wire  _GEN_219; // @[AsyncQueue.scala 113:25]
  wire  _GEN_220; // @[AsyncQueue.scala 113:25]
  wire  _GEN_221; // @[AsyncQueue.scala 113:25]
  wire  _GEN_222; // @[AsyncQueue.scala 113:25]
  wire  _GEN_223; // @[AsyncQueue.scala 113:25]
  wire  _GEN_224; // @[AsyncQueue.scala 113:25]
  wire  _GEN_225; // @[AsyncQueue.scala 113:25]
  wire  _GEN_226; // @[AsyncQueue.scala 113:25]
  wire  _GEN_227; // @[AsyncQueue.scala 113:25]
  wire  _GEN_228; // @[AsyncQueue.scala 113:25]
  wire  _GEN_229; // @[AsyncQueue.scala 113:25]
  wire  _GEN_230; // @[AsyncQueue.scala 113:25]
  wire  _GEN_231; // @[AsyncQueue.scala 113:25]
  wire  _GEN_232; // @[AsyncQueue.scala 113:25]
  wire  _GEN_233; // @[AsyncQueue.scala 113:25]
  wire  _GEN_234; // @[AsyncQueue.scala 113:25]
  wire  _GEN_235; // @[AsyncQueue.scala 113:25]
  wire  _GEN_236; // @[AsyncQueue.scala 113:25]
  wire  _GEN_237; // @[AsyncQueue.scala 113:25]
  wire  _GEN_238; // @[AsyncQueue.scala 113:25]
  wire  _GEN_239; // @[AsyncQueue.scala 113:25]
  wire  _GEN_240; // @[AsyncQueue.scala 113:25]
  wire  _GEN_241; // @[AsyncQueue.scala 113:25]
  wire  _GEN_242; // @[AsyncQueue.scala 113:25]
  wire  _GEN_243; // @[AsyncQueue.scala 113:25]
  wire  _GEN_244; // @[AsyncQueue.scala 113:25]
  wire  _GEN_245; // @[AsyncQueue.scala 113:25]
  wire  _GEN_246; // @[AsyncQueue.scala 113:25]
  wire  _GEN_247; // @[AsyncQueue.scala 113:25]
  wire  _GEN_248; // @[AsyncQueue.scala 113:25]
  wire  _GEN_249; // @[AsyncQueue.scala 113:25]
  wire  _GEN_250; // @[AsyncQueue.scala 113:25]
  wire  _GEN_251; // @[AsyncQueue.scala 113:25]
  wire  _GEN_252; // @[AsyncQueue.scala 113:25]
  wire  _GEN_253; // @[AsyncQueue.scala 113:25]
  wire  _GEN_254; // @[AsyncQueue.scala 113:25]
  wire  _GEN_255; // @[AsyncQueue.scala 113:25]
  wire  deq_bits_nxt; // @[AsyncQueue.scala 113:25]
  wire  valid_reg_1; // @[AsyncQueue.scala 116:59]
  wire  _T_293; // @[AsyncQueue.scala 117:29]
  wire  _T_298; // @[AsyncQueue.scala 127:37]
  wire  _T_299; // @[AsyncQueue.scala 127:34]
  wire  _T_318; // @[AsyncQueue.scala 139:59]
  wire  _T_291; // @[ShiftReg.scala 50:24]
  AsyncResetRegVec_w9_i0 ridx_bin ( // @[AsyncResetReg.scala 110:21]
    .clock(ridx_bin_clock),
    .reset(ridx_bin_reset),
    .io_d(ridx_bin_io_d),
    .io_q(ridx_bin_io_q),
    .io_en(ridx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w9_d3_i0 widx_gray ( // @[ShiftReg.scala 47:23]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q)
  );
  SynchronizerShiftReg_w1_d1 deq_bits_reg ( // @[ShiftReg.scala 47:23]
    .clock(deq_bits_reg_clock),
    .io_d(deq_bits_reg_io_d),
    .io_q(deq_bits_reg_io_q)
  );
  AsyncResetRegVec_w1_i0 valid_reg ( // @[AsyncResetReg.scala 110:21]
    .clock(valid_reg_clock),
    .reset(valid_reg_reset),
    .io_d(valid_reg_io_d),
    .io_q(valid_reg_io_q),
    .io_en(valid_reg_io_en)
  );
  AsyncResetRegVec_w9_i0 ridx_gray ( // @[AsyncResetReg.scala 110:21]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q),
    .io_en(ridx_gray_io_en)
  );
  AsyncValidSync_3 AsyncValidSync ( // @[AsyncQueue.scala 124:31]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_4 AsyncValidSync_1 ( // @[AsyncQueue.scala 125:31]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_5 AsyncValidSync_2 ( // @[AsyncQueue.scala 126:31]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  AsyncResetRegVec_w1_i0 AsyncResetRegVec_w1_i0 ( // @[AsyncResetReg.scala 110:21]
    .clock(AsyncResetRegVec_w1_i0_clock),
    .reset(AsyncResetRegVec_w1_i0_reset),
    .io_d(AsyncResetRegVec_w1_i0_io_d),
    .io_q(AsyncResetRegVec_w1_i0_io_q),
    .io_en(AsyncResetRegVec_w1_i0_io_en)
  );
  assign _T_272 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 30:37]
  assign source_ready = AsyncValidSync_2_io_out;
  assign _T_274 = source_ready == 1'h0; // @[AsyncQueue.scala 99:49]
  assign _GEN_256 = {{8'd0}, _T_272}; // @[AsyncQueue.scala 11:47]
  assign _T_279 = ridx_bin_io_q + _GEN_256; // @[AsyncQueue.scala 11:47]
  assign _T_280 = _T_279[8:0]; // @[AsyncQueue.scala 11:47]
  assign _T_281 = _T_274 ? 9'h0 : _T_280; // @[AsyncQueue.scala 11:23]
  assign _T_283 = _T_281 >> 1'h1; // @[AsyncQueue.scala 12:32]
  assign ridx = _T_281 ^ _T_283; // @[AsyncQueue.scala 12:17]
  assign widx = widx_gray_io_q; // @[ShiftReg.scala 50:24]
  assign _T_285 = ridx != widx; // @[AsyncQueue.scala 101:36]
  assign valid = source_ready & _T_285; // @[AsyncQueue.scala 101:28]
  assign _T_286 = ridx[7:0]; // @[AsyncQueue.scala 107:48]
  assign _T_287 = ridx[8]; // @[AsyncQueue.scala 107:67]
  assign _GEN_257 = {{7'd0}, _T_287}; // @[AsyncQueue.scala 107:80]
  assign _T_288 = _GEN_257 << 7; // @[AsyncQueue.scala 107:80]
  assign index = _T_286 ^ _T_288; // @[AsyncQueue.scala 107:60]
  assign _GEN_1 = 8'h1 == index ? io_mem_1 : io_mem_0; // @[AsyncQueue.scala 113:25]
  assign _GEN_2 = 8'h2 == index ? io_mem_2 : _GEN_1; // @[AsyncQueue.scala 113:25]
  assign _GEN_3 = 8'h3 == index ? io_mem_3 : _GEN_2; // @[AsyncQueue.scala 113:25]
  assign _GEN_4 = 8'h4 == index ? io_mem_4 : _GEN_3; // @[AsyncQueue.scala 113:25]
  assign _GEN_5 = 8'h5 == index ? io_mem_5 : _GEN_4; // @[AsyncQueue.scala 113:25]
  assign _GEN_6 = 8'h6 == index ? io_mem_6 : _GEN_5; // @[AsyncQueue.scala 113:25]
  assign _GEN_7 = 8'h7 == index ? io_mem_7 : _GEN_6; // @[AsyncQueue.scala 113:25]
  assign _GEN_8 = 8'h8 == index ? io_mem_8 : _GEN_7; // @[AsyncQueue.scala 113:25]
  assign _GEN_9 = 8'h9 == index ? io_mem_9 : _GEN_8; // @[AsyncQueue.scala 113:25]
  assign _GEN_10 = 8'ha == index ? io_mem_10 : _GEN_9; // @[AsyncQueue.scala 113:25]
  assign _GEN_11 = 8'hb == index ? io_mem_11 : _GEN_10; // @[AsyncQueue.scala 113:25]
  assign _GEN_12 = 8'hc == index ? io_mem_12 : _GEN_11; // @[AsyncQueue.scala 113:25]
  assign _GEN_13 = 8'hd == index ? io_mem_13 : _GEN_12; // @[AsyncQueue.scala 113:25]
  assign _GEN_14 = 8'he == index ? io_mem_14 : _GEN_13; // @[AsyncQueue.scala 113:25]
  assign _GEN_15 = 8'hf == index ? io_mem_15 : _GEN_14; // @[AsyncQueue.scala 113:25]
  assign _GEN_16 = 8'h10 == index ? io_mem_16 : _GEN_15; // @[AsyncQueue.scala 113:25]
  assign _GEN_17 = 8'h11 == index ? io_mem_17 : _GEN_16; // @[AsyncQueue.scala 113:25]
  assign _GEN_18 = 8'h12 == index ? io_mem_18 : _GEN_17; // @[AsyncQueue.scala 113:25]
  assign _GEN_19 = 8'h13 == index ? io_mem_19 : _GEN_18; // @[AsyncQueue.scala 113:25]
  assign _GEN_20 = 8'h14 == index ? io_mem_20 : _GEN_19; // @[AsyncQueue.scala 113:25]
  assign _GEN_21 = 8'h15 == index ? io_mem_21 : _GEN_20; // @[AsyncQueue.scala 113:25]
  assign _GEN_22 = 8'h16 == index ? io_mem_22 : _GEN_21; // @[AsyncQueue.scala 113:25]
  assign _GEN_23 = 8'h17 == index ? io_mem_23 : _GEN_22; // @[AsyncQueue.scala 113:25]
  assign _GEN_24 = 8'h18 == index ? io_mem_24 : _GEN_23; // @[AsyncQueue.scala 113:25]
  assign _GEN_25 = 8'h19 == index ? io_mem_25 : _GEN_24; // @[AsyncQueue.scala 113:25]
  assign _GEN_26 = 8'h1a == index ? io_mem_26 : _GEN_25; // @[AsyncQueue.scala 113:25]
  assign _GEN_27 = 8'h1b == index ? io_mem_27 : _GEN_26; // @[AsyncQueue.scala 113:25]
  assign _GEN_28 = 8'h1c == index ? io_mem_28 : _GEN_27; // @[AsyncQueue.scala 113:25]
  assign _GEN_29 = 8'h1d == index ? io_mem_29 : _GEN_28; // @[AsyncQueue.scala 113:25]
  assign _GEN_30 = 8'h1e == index ? io_mem_30 : _GEN_29; // @[AsyncQueue.scala 113:25]
  assign _GEN_31 = 8'h1f == index ? io_mem_31 : _GEN_30; // @[AsyncQueue.scala 113:25]
  assign _GEN_32 = 8'h20 == index ? io_mem_32 : _GEN_31; // @[AsyncQueue.scala 113:25]
  assign _GEN_33 = 8'h21 == index ? io_mem_33 : _GEN_32; // @[AsyncQueue.scala 113:25]
  assign _GEN_34 = 8'h22 == index ? io_mem_34 : _GEN_33; // @[AsyncQueue.scala 113:25]
  assign _GEN_35 = 8'h23 == index ? io_mem_35 : _GEN_34; // @[AsyncQueue.scala 113:25]
  assign _GEN_36 = 8'h24 == index ? io_mem_36 : _GEN_35; // @[AsyncQueue.scala 113:25]
  assign _GEN_37 = 8'h25 == index ? io_mem_37 : _GEN_36; // @[AsyncQueue.scala 113:25]
  assign _GEN_38 = 8'h26 == index ? io_mem_38 : _GEN_37; // @[AsyncQueue.scala 113:25]
  assign _GEN_39 = 8'h27 == index ? io_mem_39 : _GEN_38; // @[AsyncQueue.scala 113:25]
  assign _GEN_40 = 8'h28 == index ? io_mem_40 : _GEN_39; // @[AsyncQueue.scala 113:25]
  assign _GEN_41 = 8'h29 == index ? io_mem_41 : _GEN_40; // @[AsyncQueue.scala 113:25]
  assign _GEN_42 = 8'h2a == index ? io_mem_42 : _GEN_41; // @[AsyncQueue.scala 113:25]
  assign _GEN_43 = 8'h2b == index ? io_mem_43 : _GEN_42; // @[AsyncQueue.scala 113:25]
  assign _GEN_44 = 8'h2c == index ? io_mem_44 : _GEN_43; // @[AsyncQueue.scala 113:25]
  assign _GEN_45 = 8'h2d == index ? io_mem_45 : _GEN_44; // @[AsyncQueue.scala 113:25]
  assign _GEN_46 = 8'h2e == index ? io_mem_46 : _GEN_45; // @[AsyncQueue.scala 113:25]
  assign _GEN_47 = 8'h2f == index ? io_mem_47 : _GEN_46; // @[AsyncQueue.scala 113:25]
  assign _GEN_48 = 8'h30 == index ? io_mem_48 : _GEN_47; // @[AsyncQueue.scala 113:25]
  assign _GEN_49 = 8'h31 == index ? io_mem_49 : _GEN_48; // @[AsyncQueue.scala 113:25]
  assign _GEN_50 = 8'h32 == index ? io_mem_50 : _GEN_49; // @[AsyncQueue.scala 113:25]
  assign _GEN_51 = 8'h33 == index ? io_mem_51 : _GEN_50; // @[AsyncQueue.scala 113:25]
  assign _GEN_52 = 8'h34 == index ? io_mem_52 : _GEN_51; // @[AsyncQueue.scala 113:25]
  assign _GEN_53 = 8'h35 == index ? io_mem_53 : _GEN_52; // @[AsyncQueue.scala 113:25]
  assign _GEN_54 = 8'h36 == index ? io_mem_54 : _GEN_53; // @[AsyncQueue.scala 113:25]
  assign _GEN_55 = 8'h37 == index ? io_mem_55 : _GEN_54; // @[AsyncQueue.scala 113:25]
  assign _GEN_56 = 8'h38 == index ? io_mem_56 : _GEN_55; // @[AsyncQueue.scala 113:25]
  assign _GEN_57 = 8'h39 == index ? io_mem_57 : _GEN_56; // @[AsyncQueue.scala 113:25]
  assign _GEN_58 = 8'h3a == index ? io_mem_58 : _GEN_57; // @[AsyncQueue.scala 113:25]
  assign _GEN_59 = 8'h3b == index ? io_mem_59 : _GEN_58; // @[AsyncQueue.scala 113:25]
  assign _GEN_60 = 8'h3c == index ? io_mem_60 : _GEN_59; // @[AsyncQueue.scala 113:25]
  assign _GEN_61 = 8'h3d == index ? io_mem_61 : _GEN_60; // @[AsyncQueue.scala 113:25]
  assign _GEN_62 = 8'h3e == index ? io_mem_62 : _GEN_61; // @[AsyncQueue.scala 113:25]
  assign _GEN_63 = 8'h3f == index ? io_mem_63 : _GEN_62; // @[AsyncQueue.scala 113:25]
  assign _GEN_64 = 8'h40 == index ? io_mem_64 : _GEN_63; // @[AsyncQueue.scala 113:25]
  assign _GEN_65 = 8'h41 == index ? io_mem_65 : _GEN_64; // @[AsyncQueue.scala 113:25]
  assign _GEN_66 = 8'h42 == index ? io_mem_66 : _GEN_65; // @[AsyncQueue.scala 113:25]
  assign _GEN_67 = 8'h43 == index ? io_mem_67 : _GEN_66; // @[AsyncQueue.scala 113:25]
  assign _GEN_68 = 8'h44 == index ? io_mem_68 : _GEN_67; // @[AsyncQueue.scala 113:25]
  assign _GEN_69 = 8'h45 == index ? io_mem_69 : _GEN_68; // @[AsyncQueue.scala 113:25]
  assign _GEN_70 = 8'h46 == index ? io_mem_70 : _GEN_69; // @[AsyncQueue.scala 113:25]
  assign _GEN_71 = 8'h47 == index ? io_mem_71 : _GEN_70; // @[AsyncQueue.scala 113:25]
  assign _GEN_72 = 8'h48 == index ? io_mem_72 : _GEN_71; // @[AsyncQueue.scala 113:25]
  assign _GEN_73 = 8'h49 == index ? io_mem_73 : _GEN_72; // @[AsyncQueue.scala 113:25]
  assign _GEN_74 = 8'h4a == index ? io_mem_74 : _GEN_73; // @[AsyncQueue.scala 113:25]
  assign _GEN_75 = 8'h4b == index ? io_mem_75 : _GEN_74; // @[AsyncQueue.scala 113:25]
  assign _GEN_76 = 8'h4c == index ? io_mem_76 : _GEN_75; // @[AsyncQueue.scala 113:25]
  assign _GEN_77 = 8'h4d == index ? io_mem_77 : _GEN_76; // @[AsyncQueue.scala 113:25]
  assign _GEN_78 = 8'h4e == index ? io_mem_78 : _GEN_77; // @[AsyncQueue.scala 113:25]
  assign _GEN_79 = 8'h4f == index ? io_mem_79 : _GEN_78; // @[AsyncQueue.scala 113:25]
  assign _GEN_80 = 8'h50 == index ? io_mem_80 : _GEN_79; // @[AsyncQueue.scala 113:25]
  assign _GEN_81 = 8'h51 == index ? io_mem_81 : _GEN_80; // @[AsyncQueue.scala 113:25]
  assign _GEN_82 = 8'h52 == index ? io_mem_82 : _GEN_81; // @[AsyncQueue.scala 113:25]
  assign _GEN_83 = 8'h53 == index ? io_mem_83 : _GEN_82; // @[AsyncQueue.scala 113:25]
  assign _GEN_84 = 8'h54 == index ? io_mem_84 : _GEN_83; // @[AsyncQueue.scala 113:25]
  assign _GEN_85 = 8'h55 == index ? io_mem_85 : _GEN_84; // @[AsyncQueue.scala 113:25]
  assign _GEN_86 = 8'h56 == index ? io_mem_86 : _GEN_85; // @[AsyncQueue.scala 113:25]
  assign _GEN_87 = 8'h57 == index ? io_mem_87 : _GEN_86; // @[AsyncQueue.scala 113:25]
  assign _GEN_88 = 8'h58 == index ? io_mem_88 : _GEN_87; // @[AsyncQueue.scala 113:25]
  assign _GEN_89 = 8'h59 == index ? io_mem_89 : _GEN_88; // @[AsyncQueue.scala 113:25]
  assign _GEN_90 = 8'h5a == index ? io_mem_90 : _GEN_89; // @[AsyncQueue.scala 113:25]
  assign _GEN_91 = 8'h5b == index ? io_mem_91 : _GEN_90; // @[AsyncQueue.scala 113:25]
  assign _GEN_92 = 8'h5c == index ? io_mem_92 : _GEN_91; // @[AsyncQueue.scala 113:25]
  assign _GEN_93 = 8'h5d == index ? io_mem_93 : _GEN_92; // @[AsyncQueue.scala 113:25]
  assign _GEN_94 = 8'h5e == index ? io_mem_94 : _GEN_93; // @[AsyncQueue.scala 113:25]
  assign _GEN_95 = 8'h5f == index ? io_mem_95 : _GEN_94; // @[AsyncQueue.scala 113:25]
  assign _GEN_96 = 8'h60 == index ? io_mem_96 : _GEN_95; // @[AsyncQueue.scala 113:25]
  assign _GEN_97 = 8'h61 == index ? io_mem_97 : _GEN_96; // @[AsyncQueue.scala 113:25]
  assign _GEN_98 = 8'h62 == index ? io_mem_98 : _GEN_97; // @[AsyncQueue.scala 113:25]
  assign _GEN_99 = 8'h63 == index ? io_mem_99 : _GEN_98; // @[AsyncQueue.scala 113:25]
  assign _GEN_100 = 8'h64 == index ? io_mem_100 : _GEN_99; // @[AsyncQueue.scala 113:25]
  assign _GEN_101 = 8'h65 == index ? io_mem_101 : _GEN_100; // @[AsyncQueue.scala 113:25]
  assign _GEN_102 = 8'h66 == index ? io_mem_102 : _GEN_101; // @[AsyncQueue.scala 113:25]
  assign _GEN_103 = 8'h67 == index ? io_mem_103 : _GEN_102; // @[AsyncQueue.scala 113:25]
  assign _GEN_104 = 8'h68 == index ? io_mem_104 : _GEN_103; // @[AsyncQueue.scala 113:25]
  assign _GEN_105 = 8'h69 == index ? io_mem_105 : _GEN_104; // @[AsyncQueue.scala 113:25]
  assign _GEN_106 = 8'h6a == index ? io_mem_106 : _GEN_105; // @[AsyncQueue.scala 113:25]
  assign _GEN_107 = 8'h6b == index ? io_mem_107 : _GEN_106; // @[AsyncQueue.scala 113:25]
  assign _GEN_108 = 8'h6c == index ? io_mem_108 : _GEN_107; // @[AsyncQueue.scala 113:25]
  assign _GEN_109 = 8'h6d == index ? io_mem_109 : _GEN_108; // @[AsyncQueue.scala 113:25]
  assign _GEN_110 = 8'h6e == index ? io_mem_110 : _GEN_109; // @[AsyncQueue.scala 113:25]
  assign _GEN_111 = 8'h6f == index ? io_mem_111 : _GEN_110; // @[AsyncQueue.scala 113:25]
  assign _GEN_112 = 8'h70 == index ? io_mem_112 : _GEN_111; // @[AsyncQueue.scala 113:25]
  assign _GEN_113 = 8'h71 == index ? io_mem_113 : _GEN_112; // @[AsyncQueue.scala 113:25]
  assign _GEN_114 = 8'h72 == index ? io_mem_114 : _GEN_113; // @[AsyncQueue.scala 113:25]
  assign _GEN_115 = 8'h73 == index ? io_mem_115 : _GEN_114; // @[AsyncQueue.scala 113:25]
  assign _GEN_116 = 8'h74 == index ? io_mem_116 : _GEN_115; // @[AsyncQueue.scala 113:25]
  assign _GEN_117 = 8'h75 == index ? io_mem_117 : _GEN_116; // @[AsyncQueue.scala 113:25]
  assign _GEN_118 = 8'h76 == index ? io_mem_118 : _GEN_117; // @[AsyncQueue.scala 113:25]
  assign _GEN_119 = 8'h77 == index ? io_mem_119 : _GEN_118; // @[AsyncQueue.scala 113:25]
  assign _GEN_120 = 8'h78 == index ? io_mem_120 : _GEN_119; // @[AsyncQueue.scala 113:25]
  assign _GEN_121 = 8'h79 == index ? io_mem_121 : _GEN_120; // @[AsyncQueue.scala 113:25]
  assign _GEN_122 = 8'h7a == index ? io_mem_122 : _GEN_121; // @[AsyncQueue.scala 113:25]
  assign _GEN_123 = 8'h7b == index ? io_mem_123 : _GEN_122; // @[AsyncQueue.scala 113:25]
  assign _GEN_124 = 8'h7c == index ? io_mem_124 : _GEN_123; // @[AsyncQueue.scala 113:25]
  assign _GEN_125 = 8'h7d == index ? io_mem_125 : _GEN_124; // @[AsyncQueue.scala 113:25]
  assign _GEN_126 = 8'h7e == index ? io_mem_126 : _GEN_125; // @[AsyncQueue.scala 113:25]
  assign _GEN_127 = 8'h7f == index ? io_mem_127 : _GEN_126; // @[AsyncQueue.scala 113:25]
  assign _GEN_128 = 8'h80 == index ? io_mem_128 : _GEN_127; // @[AsyncQueue.scala 113:25]
  assign _GEN_129 = 8'h81 == index ? io_mem_129 : _GEN_128; // @[AsyncQueue.scala 113:25]
  assign _GEN_130 = 8'h82 == index ? io_mem_130 : _GEN_129; // @[AsyncQueue.scala 113:25]
  assign _GEN_131 = 8'h83 == index ? io_mem_131 : _GEN_130; // @[AsyncQueue.scala 113:25]
  assign _GEN_132 = 8'h84 == index ? io_mem_132 : _GEN_131; // @[AsyncQueue.scala 113:25]
  assign _GEN_133 = 8'h85 == index ? io_mem_133 : _GEN_132; // @[AsyncQueue.scala 113:25]
  assign _GEN_134 = 8'h86 == index ? io_mem_134 : _GEN_133; // @[AsyncQueue.scala 113:25]
  assign _GEN_135 = 8'h87 == index ? io_mem_135 : _GEN_134; // @[AsyncQueue.scala 113:25]
  assign _GEN_136 = 8'h88 == index ? io_mem_136 : _GEN_135; // @[AsyncQueue.scala 113:25]
  assign _GEN_137 = 8'h89 == index ? io_mem_137 : _GEN_136; // @[AsyncQueue.scala 113:25]
  assign _GEN_138 = 8'h8a == index ? io_mem_138 : _GEN_137; // @[AsyncQueue.scala 113:25]
  assign _GEN_139 = 8'h8b == index ? io_mem_139 : _GEN_138; // @[AsyncQueue.scala 113:25]
  assign _GEN_140 = 8'h8c == index ? io_mem_140 : _GEN_139; // @[AsyncQueue.scala 113:25]
  assign _GEN_141 = 8'h8d == index ? io_mem_141 : _GEN_140; // @[AsyncQueue.scala 113:25]
  assign _GEN_142 = 8'h8e == index ? io_mem_142 : _GEN_141; // @[AsyncQueue.scala 113:25]
  assign _GEN_143 = 8'h8f == index ? io_mem_143 : _GEN_142; // @[AsyncQueue.scala 113:25]
  assign _GEN_144 = 8'h90 == index ? io_mem_144 : _GEN_143; // @[AsyncQueue.scala 113:25]
  assign _GEN_145 = 8'h91 == index ? io_mem_145 : _GEN_144; // @[AsyncQueue.scala 113:25]
  assign _GEN_146 = 8'h92 == index ? io_mem_146 : _GEN_145; // @[AsyncQueue.scala 113:25]
  assign _GEN_147 = 8'h93 == index ? io_mem_147 : _GEN_146; // @[AsyncQueue.scala 113:25]
  assign _GEN_148 = 8'h94 == index ? io_mem_148 : _GEN_147; // @[AsyncQueue.scala 113:25]
  assign _GEN_149 = 8'h95 == index ? io_mem_149 : _GEN_148; // @[AsyncQueue.scala 113:25]
  assign _GEN_150 = 8'h96 == index ? io_mem_150 : _GEN_149; // @[AsyncQueue.scala 113:25]
  assign _GEN_151 = 8'h97 == index ? io_mem_151 : _GEN_150; // @[AsyncQueue.scala 113:25]
  assign _GEN_152 = 8'h98 == index ? io_mem_152 : _GEN_151; // @[AsyncQueue.scala 113:25]
  assign _GEN_153 = 8'h99 == index ? io_mem_153 : _GEN_152; // @[AsyncQueue.scala 113:25]
  assign _GEN_154 = 8'h9a == index ? io_mem_154 : _GEN_153; // @[AsyncQueue.scala 113:25]
  assign _GEN_155 = 8'h9b == index ? io_mem_155 : _GEN_154; // @[AsyncQueue.scala 113:25]
  assign _GEN_156 = 8'h9c == index ? io_mem_156 : _GEN_155; // @[AsyncQueue.scala 113:25]
  assign _GEN_157 = 8'h9d == index ? io_mem_157 : _GEN_156; // @[AsyncQueue.scala 113:25]
  assign _GEN_158 = 8'h9e == index ? io_mem_158 : _GEN_157; // @[AsyncQueue.scala 113:25]
  assign _GEN_159 = 8'h9f == index ? io_mem_159 : _GEN_158; // @[AsyncQueue.scala 113:25]
  assign _GEN_160 = 8'ha0 == index ? io_mem_160 : _GEN_159; // @[AsyncQueue.scala 113:25]
  assign _GEN_161 = 8'ha1 == index ? io_mem_161 : _GEN_160; // @[AsyncQueue.scala 113:25]
  assign _GEN_162 = 8'ha2 == index ? io_mem_162 : _GEN_161; // @[AsyncQueue.scala 113:25]
  assign _GEN_163 = 8'ha3 == index ? io_mem_163 : _GEN_162; // @[AsyncQueue.scala 113:25]
  assign _GEN_164 = 8'ha4 == index ? io_mem_164 : _GEN_163; // @[AsyncQueue.scala 113:25]
  assign _GEN_165 = 8'ha5 == index ? io_mem_165 : _GEN_164; // @[AsyncQueue.scala 113:25]
  assign _GEN_166 = 8'ha6 == index ? io_mem_166 : _GEN_165; // @[AsyncQueue.scala 113:25]
  assign _GEN_167 = 8'ha7 == index ? io_mem_167 : _GEN_166; // @[AsyncQueue.scala 113:25]
  assign _GEN_168 = 8'ha8 == index ? io_mem_168 : _GEN_167; // @[AsyncQueue.scala 113:25]
  assign _GEN_169 = 8'ha9 == index ? io_mem_169 : _GEN_168; // @[AsyncQueue.scala 113:25]
  assign _GEN_170 = 8'haa == index ? io_mem_170 : _GEN_169; // @[AsyncQueue.scala 113:25]
  assign _GEN_171 = 8'hab == index ? io_mem_171 : _GEN_170; // @[AsyncQueue.scala 113:25]
  assign _GEN_172 = 8'hac == index ? io_mem_172 : _GEN_171; // @[AsyncQueue.scala 113:25]
  assign _GEN_173 = 8'had == index ? io_mem_173 : _GEN_172; // @[AsyncQueue.scala 113:25]
  assign _GEN_174 = 8'hae == index ? io_mem_174 : _GEN_173; // @[AsyncQueue.scala 113:25]
  assign _GEN_175 = 8'haf == index ? io_mem_175 : _GEN_174; // @[AsyncQueue.scala 113:25]
  assign _GEN_176 = 8'hb0 == index ? io_mem_176 : _GEN_175; // @[AsyncQueue.scala 113:25]
  assign _GEN_177 = 8'hb1 == index ? io_mem_177 : _GEN_176; // @[AsyncQueue.scala 113:25]
  assign _GEN_178 = 8'hb2 == index ? io_mem_178 : _GEN_177; // @[AsyncQueue.scala 113:25]
  assign _GEN_179 = 8'hb3 == index ? io_mem_179 : _GEN_178; // @[AsyncQueue.scala 113:25]
  assign _GEN_180 = 8'hb4 == index ? io_mem_180 : _GEN_179; // @[AsyncQueue.scala 113:25]
  assign _GEN_181 = 8'hb5 == index ? io_mem_181 : _GEN_180; // @[AsyncQueue.scala 113:25]
  assign _GEN_182 = 8'hb6 == index ? io_mem_182 : _GEN_181; // @[AsyncQueue.scala 113:25]
  assign _GEN_183 = 8'hb7 == index ? io_mem_183 : _GEN_182; // @[AsyncQueue.scala 113:25]
  assign _GEN_184 = 8'hb8 == index ? io_mem_184 : _GEN_183; // @[AsyncQueue.scala 113:25]
  assign _GEN_185 = 8'hb9 == index ? io_mem_185 : _GEN_184; // @[AsyncQueue.scala 113:25]
  assign _GEN_186 = 8'hba == index ? io_mem_186 : _GEN_185; // @[AsyncQueue.scala 113:25]
  assign _GEN_187 = 8'hbb == index ? io_mem_187 : _GEN_186; // @[AsyncQueue.scala 113:25]
  assign _GEN_188 = 8'hbc == index ? io_mem_188 : _GEN_187; // @[AsyncQueue.scala 113:25]
  assign _GEN_189 = 8'hbd == index ? io_mem_189 : _GEN_188; // @[AsyncQueue.scala 113:25]
  assign _GEN_190 = 8'hbe == index ? io_mem_190 : _GEN_189; // @[AsyncQueue.scala 113:25]
  assign _GEN_191 = 8'hbf == index ? io_mem_191 : _GEN_190; // @[AsyncQueue.scala 113:25]
  assign _GEN_192 = 8'hc0 == index ? io_mem_192 : _GEN_191; // @[AsyncQueue.scala 113:25]
  assign _GEN_193 = 8'hc1 == index ? io_mem_193 : _GEN_192; // @[AsyncQueue.scala 113:25]
  assign _GEN_194 = 8'hc2 == index ? io_mem_194 : _GEN_193; // @[AsyncQueue.scala 113:25]
  assign _GEN_195 = 8'hc3 == index ? io_mem_195 : _GEN_194; // @[AsyncQueue.scala 113:25]
  assign _GEN_196 = 8'hc4 == index ? io_mem_196 : _GEN_195; // @[AsyncQueue.scala 113:25]
  assign _GEN_197 = 8'hc5 == index ? io_mem_197 : _GEN_196; // @[AsyncQueue.scala 113:25]
  assign _GEN_198 = 8'hc6 == index ? io_mem_198 : _GEN_197; // @[AsyncQueue.scala 113:25]
  assign _GEN_199 = 8'hc7 == index ? io_mem_199 : _GEN_198; // @[AsyncQueue.scala 113:25]
  assign _GEN_200 = 8'hc8 == index ? io_mem_200 : _GEN_199; // @[AsyncQueue.scala 113:25]
  assign _GEN_201 = 8'hc9 == index ? io_mem_201 : _GEN_200; // @[AsyncQueue.scala 113:25]
  assign _GEN_202 = 8'hca == index ? io_mem_202 : _GEN_201; // @[AsyncQueue.scala 113:25]
  assign _GEN_203 = 8'hcb == index ? io_mem_203 : _GEN_202; // @[AsyncQueue.scala 113:25]
  assign _GEN_204 = 8'hcc == index ? io_mem_204 : _GEN_203; // @[AsyncQueue.scala 113:25]
  assign _GEN_205 = 8'hcd == index ? io_mem_205 : _GEN_204; // @[AsyncQueue.scala 113:25]
  assign _GEN_206 = 8'hce == index ? io_mem_206 : _GEN_205; // @[AsyncQueue.scala 113:25]
  assign _GEN_207 = 8'hcf == index ? io_mem_207 : _GEN_206; // @[AsyncQueue.scala 113:25]
  assign _GEN_208 = 8'hd0 == index ? io_mem_208 : _GEN_207; // @[AsyncQueue.scala 113:25]
  assign _GEN_209 = 8'hd1 == index ? io_mem_209 : _GEN_208; // @[AsyncQueue.scala 113:25]
  assign _GEN_210 = 8'hd2 == index ? io_mem_210 : _GEN_209; // @[AsyncQueue.scala 113:25]
  assign _GEN_211 = 8'hd3 == index ? io_mem_211 : _GEN_210; // @[AsyncQueue.scala 113:25]
  assign _GEN_212 = 8'hd4 == index ? io_mem_212 : _GEN_211; // @[AsyncQueue.scala 113:25]
  assign _GEN_213 = 8'hd5 == index ? io_mem_213 : _GEN_212; // @[AsyncQueue.scala 113:25]
  assign _GEN_214 = 8'hd6 == index ? io_mem_214 : _GEN_213; // @[AsyncQueue.scala 113:25]
  assign _GEN_215 = 8'hd7 == index ? io_mem_215 : _GEN_214; // @[AsyncQueue.scala 113:25]
  assign _GEN_216 = 8'hd8 == index ? io_mem_216 : _GEN_215; // @[AsyncQueue.scala 113:25]
  assign _GEN_217 = 8'hd9 == index ? io_mem_217 : _GEN_216; // @[AsyncQueue.scala 113:25]
  assign _GEN_218 = 8'hda == index ? io_mem_218 : _GEN_217; // @[AsyncQueue.scala 113:25]
  assign _GEN_219 = 8'hdb == index ? io_mem_219 : _GEN_218; // @[AsyncQueue.scala 113:25]
  assign _GEN_220 = 8'hdc == index ? io_mem_220 : _GEN_219; // @[AsyncQueue.scala 113:25]
  assign _GEN_221 = 8'hdd == index ? io_mem_221 : _GEN_220; // @[AsyncQueue.scala 113:25]
  assign _GEN_222 = 8'hde == index ? io_mem_222 : _GEN_221; // @[AsyncQueue.scala 113:25]
  assign _GEN_223 = 8'hdf == index ? io_mem_223 : _GEN_222; // @[AsyncQueue.scala 113:25]
  assign _GEN_224 = 8'he0 == index ? io_mem_224 : _GEN_223; // @[AsyncQueue.scala 113:25]
  assign _GEN_225 = 8'he1 == index ? io_mem_225 : _GEN_224; // @[AsyncQueue.scala 113:25]
  assign _GEN_226 = 8'he2 == index ? io_mem_226 : _GEN_225; // @[AsyncQueue.scala 113:25]
  assign _GEN_227 = 8'he3 == index ? io_mem_227 : _GEN_226; // @[AsyncQueue.scala 113:25]
  assign _GEN_228 = 8'he4 == index ? io_mem_228 : _GEN_227; // @[AsyncQueue.scala 113:25]
  assign _GEN_229 = 8'he5 == index ? io_mem_229 : _GEN_228; // @[AsyncQueue.scala 113:25]
  assign _GEN_230 = 8'he6 == index ? io_mem_230 : _GEN_229; // @[AsyncQueue.scala 113:25]
  assign _GEN_231 = 8'he7 == index ? io_mem_231 : _GEN_230; // @[AsyncQueue.scala 113:25]
  assign _GEN_232 = 8'he8 == index ? io_mem_232 : _GEN_231; // @[AsyncQueue.scala 113:25]
  assign _GEN_233 = 8'he9 == index ? io_mem_233 : _GEN_232; // @[AsyncQueue.scala 113:25]
  assign _GEN_234 = 8'hea == index ? io_mem_234 : _GEN_233; // @[AsyncQueue.scala 113:25]
  assign _GEN_235 = 8'heb == index ? io_mem_235 : _GEN_234; // @[AsyncQueue.scala 113:25]
  assign _GEN_236 = 8'hec == index ? io_mem_236 : _GEN_235; // @[AsyncQueue.scala 113:25]
  assign _GEN_237 = 8'hed == index ? io_mem_237 : _GEN_236; // @[AsyncQueue.scala 113:25]
  assign _GEN_238 = 8'hee == index ? io_mem_238 : _GEN_237; // @[AsyncQueue.scala 113:25]
  assign _GEN_239 = 8'hef == index ? io_mem_239 : _GEN_238; // @[AsyncQueue.scala 113:25]
  assign _GEN_240 = 8'hf0 == index ? io_mem_240 : _GEN_239; // @[AsyncQueue.scala 113:25]
  assign _GEN_241 = 8'hf1 == index ? io_mem_241 : _GEN_240; // @[AsyncQueue.scala 113:25]
  assign _GEN_242 = 8'hf2 == index ? io_mem_242 : _GEN_241; // @[AsyncQueue.scala 113:25]
  assign _GEN_243 = 8'hf3 == index ? io_mem_243 : _GEN_242; // @[AsyncQueue.scala 113:25]
  assign _GEN_244 = 8'hf4 == index ? io_mem_244 : _GEN_243; // @[AsyncQueue.scala 113:25]
  assign _GEN_245 = 8'hf5 == index ? io_mem_245 : _GEN_244; // @[AsyncQueue.scala 113:25]
  assign _GEN_246 = 8'hf6 == index ? io_mem_246 : _GEN_245; // @[AsyncQueue.scala 113:25]
  assign _GEN_247 = 8'hf7 == index ? io_mem_247 : _GEN_246; // @[AsyncQueue.scala 113:25]
  assign _GEN_248 = 8'hf8 == index ? io_mem_248 : _GEN_247; // @[AsyncQueue.scala 113:25]
  assign _GEN_249 = 8'hf9 == index ? io_mem_249 : _GEN_248; // @[AsyncQueue.scala 113:25]
  assign _GEN_250 = 8'hfa == index ? io_mem_250 : _GEN_249; // @[AsyncQueue.scala 113:25]
  assign _GEN_251 = 8'hfb == index ? io_mem_251 : _GEN_250; // @[AsyncQueue.scala 113:25]
  assign _GEN_252 = 8'hfc == index ? io_mem_252 : _GEN_251; // @[AsyncQueue.scala 113:25]
  assign _GEN_253 = 8'hfd == index ? io_mem_253 : _GEN_252; // @[AsyncQueue.scala 113:25]
  assign _GEN_254 = 8'hfe == index ? io_mem_254 : _GEN_253; // @[AsyncQueue.scala 113:25]
  assign _GEN_255 = 8'hff == index ? io_mem_255 : _GEN_254; // @[AsyncQueue.scala 113:25]
  assign deq_bits_nxt = valid ? _GEN_255 : io_deq_bits; // @[AsyncQueue.scala 113:25]
  assign valid_reg_1 = valid_reg_io_q; // @[AsyncQueue.scala 116:59]
  assign _T_293 = valid_reg_1 & source_ready; // @[AsyncQueue.scala 117:29]
  assign _T_298 = io_source_reset_n == 1'h0; // @[AsyncQueue.scala 127:37]
  assign _T_299 = reset | _T_298; // @[AsyncQueue.scala 127:34]
  assign _T_318 = io_widx == io_ridx; // @[AsyncQueue.scala 139:59]
  assign _T_291 = deq_bits_reg_io_q; // @[ShiftReg.scala 50:24]
  assign io_deq_valid = _T_293;
  assign io_deq_bits = _T_291;
  assign io_ridx = ridx_gray_io_q;
  assign io_ridx_valid = AsyncValidSync_io_out;
  assign ridx_bin_clock = clock;
  assign ridx_bin_reset = reset;
  assign ridx_bin_io_d = _T_281;
  assign ridx_bin_io_en = 1'h1;
  assign widx_gray_clock = clock;
  assign widx_gray_reset = reset;
  assign widx_gray_io_d = io_widx;
  assign deq_bits_reg_clock = clock;
  assign deq_bits_reg_io_d = deq_bits_nxt;
  assign valid_reg_clock = clock;
  assign valid_reg_reset = reset;
  assign valid_reg_io_d = valid;
  assign valid_reg_io_en = 1'h1;
  assign ridx_gray_clock = clock;
  assign ridx_gray_reset = reset;
  assign ridx_gray_io_d = ridx;
  assign ridx_gray_io_en = 1'h1;
  assign AsyncValidSync_clock = clock;
  assign AsyncValidSync_reset = _T_299;
  assign AsyncValidSync_1_clock = clock;
  assign AsyncValidSync_1_reset = _T_299;
  assign AsyncValidSync_1_io_in = io_widx_valid;
  assign AsyncValidSync_2_clock = clock;
  assign AsyncValidSync_2_reset = reset;
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out;
  assign AsyncResetRegVec_w1_i0_clock = clock;
  assign AsyncResetRegVec_w1_i0_reset = reset;
  assign AsyncResetRegVec_w1_i0_io_d = _T_318;
  assign AsyncResetRegVec_w1_i0_io_en = 1'h1;
endmodule
module AsyncQueue(
  input   io_enq_clock,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits,
  input   io_deq_clock,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits
);
  wire  source_clock; // @[AsyncQueue.scala 155:22]
  wire  source_reset; // @[AsyncQueue.scala 155:22]
  wire  source_io_enq_ready; // @[AsyncQueue.scala 155:22]
  wire  source_io_enq_valid; // @[AsyncQueue.scala 155:22]
  wire  source_io_enq_bits; // @[AsyncQueue.scala 155:22]
  wire [8:0] source_io_ridx; // @[AsyncQueue.scala 155:22]
  wire [8:0] source_io_widx; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_0; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_1; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_2; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_3; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_4; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_5; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_6; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_7; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_8; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_9; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_10; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_11; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_12; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_13; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_14; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_15; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_16; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_17; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_18; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_19; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_20; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_21; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_22; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_23; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_24; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_25; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_26; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_27; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_28; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_29; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_30; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_31; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_32; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_33; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_34; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_35; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_36; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_37; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_38; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_39; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_40; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_41; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_42; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_43; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_44; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_45; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_46; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_47; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_48; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_49; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_50; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_51; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_52; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_53; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_54; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_55; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_56; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_57; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_58; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_59; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_60; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_61; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_62; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_63; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_64; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_65; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_66; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_67; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_68; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_69; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_70; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_71; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_72; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_73; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_74; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_75; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_76; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_77; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_78; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_79; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_80; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_81; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_82; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_83; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_84; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_85; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_86; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_87; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_88; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_89; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_90; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_91; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_92; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_93; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_94; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_95; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_96; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_97; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_98; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_99; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_100; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_101; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_102; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_103; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_104; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_105; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_106; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_107; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_108; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_109; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_110; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_111; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_112; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_113; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_114; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_115; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_116; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_117; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_118; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_119; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_120; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_121; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_122; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_123; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_124; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_125; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_126; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_127; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_128; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_129; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_130; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_131; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_132; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_133; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_134; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_135; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_136; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_137; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_138; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_139; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_140; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_141; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_142; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_143; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_144; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_145; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_146; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_147; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_148; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_149; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_150; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_151; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_152; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_153; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_154; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_155; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_156; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_157; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_158; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_159; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_160; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_161; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_162; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_163; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_164; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_165; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_166; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_167; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_168; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_169; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_170; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_171; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_172; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_173; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_174; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_175; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_176; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_177; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_178; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_179; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_180; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_181; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_182; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_183; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_184; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_185; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_186; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_187; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_188; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_189; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_190; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_191; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_192; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_193; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_194; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_195; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_196; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_197; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_198; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_199; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_200; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_201; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_202; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_203; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_204; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_205; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_206; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_207; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_208; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_209; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_210; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_211; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_212; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_213; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_214; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_215; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_216; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_217; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_218; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_219; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_220; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_221; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_222; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_223; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_224; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_225; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_226; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_227; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_228; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_229; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_230; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_231; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_232; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_233; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_234; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_235; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_236; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_237; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_238; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_239; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_240; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_241; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_242; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_243; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_244; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_245; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_246; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_247; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_248; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_249; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_250; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_251; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_252; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_253; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_254; // @[AsyncQueue.scala 155:22]
  wire  source_io_mem_255; // @[AsyncQueue.scala 155:22]
  wire  source_io_sink_reset_n; // @[AsyncQueue.scala 155:22]
  wire  source_io_ridx_valid; // @[AsyncQueue.scala 155:22]
  wire  source_io_widx_valid; // @[AsyncQueue.scala 155:22]
  wire  sink_clock; // @[AsyncQueue.scala 156:22]
  wire  sink_reset; // @[AsyncQueue.scala 156:22]
  wire  sink_io_deq_ready; // @[AsyncQueue.scala 156:22]
  wire  sink_io_deq_valid; // @[AsyncQueue.scala 156:22]
  wire  sink_io_deq_bits; // @[AsyncQueue.scala 156:22]
  wire [8:0] sink_io_ridx; // @[AsyncQueue.scala 156:22]
  wire [8:0] sink_io_widx; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_0; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_1; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_2; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_3; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_4; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_5; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_6; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_7; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_8; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_9; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_10; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_11; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_12; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_13; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_14; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_15; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_16; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_17; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_18; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_19; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_20; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_21; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_22; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_23; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_24; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_25; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_26; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_27; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_28; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_29; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_30; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_31; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_32; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_33; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_34; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_35; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_36; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_37; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_38; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_39; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_40; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_41; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_42; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_43; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_44; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_45; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_46; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_47; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_48; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_49; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_50; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_51; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_52; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_53; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_54; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_55; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_56; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_57; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_58; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_59; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_60; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_61; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_62; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_63; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_64; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_65; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_66; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_67; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_68; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_69; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_70; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_71; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_72; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_73; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_74; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_75; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_76; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_77; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_78; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_79; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_80; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_81; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_82; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_83; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_84; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_85; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_86; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_87; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_88; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_89; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_90; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_91; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_92; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_93; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_94; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_95; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_96; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_97; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_98; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_99; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_100; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_101; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_102; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_103; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_104; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_105; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_106; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_107; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_108; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_109; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_110; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_111; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_112; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_113; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_114; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_115; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_116; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_117; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_118; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_119; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_120; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_121; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_122; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_123; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_124; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_125; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_126; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_127; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_128; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_129; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_130; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_131; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_132; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_133; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_134; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_135; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_136; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_137; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_138; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_139; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_140; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_141; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_142; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_143; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_144; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_145; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_146; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_147; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_148; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_149; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_150; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_151; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_152; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_153; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_154; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_155; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_156; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_157; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_158; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_159; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_160; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_161; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_162; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_163; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_164; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_165; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_166; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_167; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_168; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_169; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_170; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_171; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_172; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_173; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_174; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_175; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_176; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_177; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_178; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_179; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_180; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_181; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_182; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_183; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_184; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_185; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_186; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_187; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_188; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_189; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_190; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_191; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_192; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_193; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_194; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_195; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_196; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_197; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_198; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_199; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_200; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_201; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_202; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_203; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_204; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_205; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_206; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_207; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_208; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_209; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_210; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_211; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_212; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_213; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_214; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_215; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_216; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_217; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_218; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_219; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_220; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_221; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_222; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_223; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_224; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_225; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_226; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_227; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_228; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_229; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_230; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_231; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_232; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_233; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_234; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_235; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_236; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_237; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_238; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_239; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_240; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_241; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_242; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_243; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_244; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_245; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_246; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_247; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_248; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_249; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_250; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_251; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_252; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_253; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_254; // @[AsyncQueue.scala 156:22]
  wire  sink_io_mem_255; // @[AsyncQueue.scala 156:22]
  wire  sink_io_source_reset_n; // @[AsyncQueue.scala 156:22]
  wire  sink_io_ridx_valid; // @[AsyncQueue.scala 156:22]
  wire  sink_io_widx_valid; // @[AsyncQueue.scala 156:22]
  AsyncQueueSource source ( // @[AsyncQueue.scala 155:22]
    .clock(source_clock),
    .reset(source_reset),
    .io_enq_ready(source_io_enq_ready),
    .io_enq_valid(source_io_enq_valid),
    .io_enq_bits(source_io_enq_bits),
    .io_ridx(source_io_ridx),
    .io_widx(source_io_widx),
    .io_mem_0(source_io_mem_0),
    .io_mem_1(source_io_mem_1),
    .io_mem_2(source_io_mem_2),
    .io_mem_3(source_io_mem_3),
    .io_mem_4(source_io_mem_4),
    .io_mem_5(source_io_mem_5),
    .io_mem_6(source_io_mem_6),
    .io_mem_7(source_io_mem_7),
    .io_mem_8(source_io_mem_8),
    .io_mem_9(source_io_mem_9),
    .io_mem_10(source_io_mem_10),
    .io_mem_11(source_io_mem_11),
    .io_mem_12(source_io_mem_12),
    .io_mem_13(source_io_mem_13),
    .io_mem_14(source_io_mem_14),
    .io_mem_15(source_io_mem_15),
    .io_mem_16(source_io_mem_16),
    .io_mem_17(source_io_mem_17),
    .io_mem_18(source_io_mem_18),
    .io_mem_19(source_io_mem_19),
    .io_mem_20(source_io_mem_20),
    .io_mem_21(source_io_mem_21),
    .io_mem_22(source_io_mem_22),
    .io_mem_23(source_io_mem_23),
    .io_mem_24(source_io_mem_24),
    .io_mem_25(source_io_mem_25),
    .io_mem_26(source_io_mem_26),
    .io_mem_27(source_io_mem_27),
    .io_mem_28(source_io_mem_28),
    .io_mem_29(source_io_mem_29),
    .io_mem_30(source_io_mem_30),
    .io_mem_31(source_io_mem_31),
    .io_mem_32(source_io_mem_32),
    .io_mem_33(source_io_mem_33),
    .io_mem_34(source_io_mem_34),
    .io_mem_35(source_io_mem_35),
    .io_mem_36(source_io_mem_36),
    .io_mem_37(source_io_mem_37),
    .io_mem_38(source_io_mem_38),
    .io_mem_39(source_io_mem_39),
    .io_mem_40(source_io_mem_40),
    .io_mem_41(source_io_mem_41),
    .io_mem_42(source_io_mem_42),
    .io_mem_43(source_io_mem_43),
    .io_mem_44(source_io_mem_44),
    .io_mem_45(source_io_mem_45),
    .io_mem_46(source_io_mem_46),
    .io_mem_47(source_io_mem_47),
    .io_mem_48(source_io_mem_48),
    .io_mem_49(source_io_mem_49),
    .io_mem_50(source_io_mem_50),
    .io_mem_51(source_io_mem_51),
    .io_mem_52(source_io_mem_52),
    .io_mem_53(source_io_mem_53),
    .io_mem_54(source_io_mem_54),
    .io_mem_55(source_io_mem_55),
    .io_mem_56(source_io_mem_56),
    .io_mem_57(source_io_mem_57),
    .io_mem_58(source_io_mem_58),
    .io_mem_59(source_io_mem_59),
    .io_mem_60(source_io_mem_60),
    .io_mem_61(source_io_mem_61),
    .io_mem_62(source_io_mem_62),
    .io_mem_63(source_io_mem_63),
    .io_mem_64(source_io_mem_64),
    .io_mem_65(source_io_mem_65),
    .io_mem_66(source_io_mem_66),
    .io_mem_67(source_io_mem_67),
    .io_mem_68(source_io_mem_68),
    .io_mem_69(source_io_mem_69),
    .io_mem_70(source_io_mem_70),
    .io_mem_71(source_io_mem_71),
    .io_mem_72(source_io_mem_72),
    .io_mem_73(source_io_mem_73),
    .io_mem_74(source_io_mem_74),
    .io_mem_75(source_io_mem_75),
    .io_mem_76(source_io_mem_76),
    .io_mem_77(source_io_mem_77),
    .io_mem_78(source_io_mem_78),
    .io_mem_79(source_io_mem_79),
    .io_mem_80(source_io_mem_80),
    .io_mem_81(source_io_mem_81),
    .io_mem_82(source_io_mem_82),
    .io_mem_83(source_io_mem_83),
    .io_mem_84(source_io_mem_84),
    .io_mem_85(source_io_mem_85),
    .io_mem_86(source_io_mem_86),
    .io_mem_87(source_io_mem_87),
    .io_mem_88(source_io_mem_88),
    .io_mem_89(source_io_mem_89),
    .io_mem_90(source_io_mem_90),
    .io_mem_91(source_io_mem_91),
    .io_mem_92(source_io_mem_92),
    .io_mem_93(source_io_mem_93),
    .io_mem_94(source_io_mem_94),
    .io_mem_95(source_io_mem_95),
    .io_mem_96(source_io_mem_96),
    .io_mem_97(source_io_mem_97),
    .io_mem_98(source_io_mem_98),
    .io_mem_99(source_io_mem_99),
    .io_mem_100(source_io_mem_100),
    .io_mem_101(source_io_mem_101),
    .io_mem_102(source_io_mem_102),
    .io_mem_103(source_io_mem_103),
    .io_mem_104(source_io_mem_104),
    .io_mem_105(source_io_mem_105),
    .io_mem_106(source_io_mem_106),
    .io_mem_107(source_io_mem_107),
    .io_mem_108(source_io_mem_108),
    .io_mem_109(source_io_mem_109),
    .io_mem_110(source_io_mem_110),
    .io_mem_111(source_io_mem_111),
    .io_mem_112(source_io_mem_112),
    .io_mem_113(source_io_mem_113),
    .io_mem_114(source_io_mem_114),
    .io_mem_115(source_io_mem_115),
    .io_mem_116(source_io_mem_116),
    .io_mem_117(source_io_mem_117),
    .io_mem_118(source_io_mem_118),
    .io_mem_119(source_io_mem_119),
    .io_mem_120(source_io_mem_120),
    .io_mem_121(source_io_mem_121),
    .io_mem_122(source_io_mem_122),
    .io_mem_123(source_io_mem_123),
    .io_mem_124(source_io_mem_124),
    .io_mem_125(source_io_mem_125),
    .io_mem_126(source_io_mem_126),
    .io_mem_127(source_io_mem_127),
    .io_mem_128(source_io_mem_128),
    .io_mem_129(source_io_mem_129),
    .io_mem_130(source_io_mem_130),
    .io_mem_131(source_io_mem_131),
    .io_mem_132(source_io_mem_132),
    .io_mem_133(source_io_mem_133),
    .io_mem_134(source_io_mem_134),
    .io_mem_135(source_io_mem_135),
    .io_mem_136(source_io_mem_136),
    .io_mem_137(source_io_mem_137),
    .io_mem_138(source_io_mem_138),
    .io_mem_139(source_io_mem_139),
    .io_mem_140(source_io_mem_140),
    .io_mem_141(source_io_mem_141),
    .io_mem_142(source_io_mem_142),
    .io_mem_143(source_io_mem_143),
    .io_mem_144(source_io_mem_144),
    .io_mem_145(source_io_mem_145),
    .io_mem_146(source_io_mem_146),
    .io_mem_147(source_io_mem_147),
    .io_mem_148(source_io_mem_148),
    .io_mem_149(source_io_mem_149),
    .io_mem_150(source_io_mem_150),
    .io_mem_151(source_io_mem_151),
    .io_mem_152(source_io_mem_152),
    .io_mem_153(source_io_mem_153),
    .io_mem_154(source_io_mem_154),
    .io_mem_155(source_io_mem_155),
    .io_mem_156(source_io_mem_156),
    .io_mem_157(source_io_mem_157),
    .io_mem_158(source_io_mem_158),
    .io_mem_159(source_io_mem_159),
    .io_mem_160(source_io_mem_160),
    .io_mem_161(source_io_mem_161),
    .io_mem_162(source_io_mem_162),
    .io_mem_163(source_io_mem_163),
    .io_mem_164(source_io_mem_164),
    .io_mem_165(source_io_mem_165),
    .io_mem_166(source_io_mem_166),
    .io_mem_167(source_io_mem_167),
    .io_mem_168(source_io_mem_168),
    .io_mem_169(source_io_mem_169),
    .io_mem_170(source_io_mem_170),
    .io_mem_171(source_io_mem_171),
    .io_mem_172(source_io_mem_172),
    .io_mem_173(source_io_mem_173),
    .io_mem_174(source_io_mem_174),
    .io_mem_175(source_io_mem_175),
    .io_mem_176(source_io_mem_176),
    .io_mem_177(source_io_mem_177),
    .io_mem_178(source_io_mem_178),
    .io_mem_179(source_io_mem_179),
    .io_mem_180(source_io_mem_180),
    .io_mem_181(source_io_mem_181),
    .io_mem_182(source_io_mem_182),
    .io_mem_183(source_io_mem_183),
    .io_mem_184(source_io_mem_184),
    .io_mem_185(source_io_mem_185),
    .io_mem_186(source_io_mem_186),
    .io_mem_187(source_io_mem_187),
    .io_mem_188(source_io_mem_188),
    .io_mem_189(source_io_mem_189),
    .io_mem_190(source_io_mem_190),
    .io_mem_191(source_io_mem_191),
    .io_mem_192(source_io_mem_192),
    .io_mem_193(source_io_mem_193),
    .io_mem_194(source_io_mem_194),
    .io_mem_195(source_io_mem_195),
    .io_mem_196(source_io_mem_196),
    .io_mem_197(source_io_mem_197),
    .io_mem_198(source_io_mem_198),
    .io_mem_199(source_io_mem_199),
    .io_mem_200(source_io_mem_200),
    .io_mem_201(source_io_mem_201),
    .io_mem_202(source_io_mem_202),
    .io_mem_203(source_io_mem_203),
    .io_mem_204(source_io_mem_204),
    .io_mem_205(source_io_mem_205),
    .io_mem_206(source_io_mem_206),
    .io_mem_207(source_io_mem_207),
    .io_mem_208(source_io_mem_208),
    .io_mem_209(source_io_mem_209),
    .io_mem_210(source_io_mem_210),
    .io_mem_211(source_io_mem_211),
    .io_mem_212(source_io_mem_212),
    .io_mem_213(source_io_mem_213),
    .io_mem_214(source_io_mem_214),
    .io_mem_215(source_io_mem_215),
    .io_mem_216(source_io_mem_216),
    .io_mem_217(source_io_mem_217),
    .io_mem_218(source_io_mem_218),
    .io_mem_219(source_io_mem_219),
    .io_mem_220(source_io_mem_220),
    .io_mem_221(source_io_mem_221),
    .io_mem_222(source_io_mem_222),
    .io_mem_223(source_io_mem_223),
    .io_mem_224(source_io_mem_224),
    .io_mem_225(source_io_mem_225),
    .io_mem_226(source_io_mem_226),
    .io_mem_227(source_io_mem_227),
    .io_mem_228(source_io_mem_228),
    .io_mem_229(source_io_mem_229),
    .io_mem_230(source_io_mem_230),
    .io_mem_231(source_io_mem_231),
    .io_mem_232(source_io_mem_232),
    .io_mem_233(source_io_mem_233),
    .io_mem_234(source_io_mem_234),
    .io_mem_235(source_io_mem_235),
    .io_mem_236(source_io_mem_236),
    .io_mem_237(source_io_mem_237),
    .io_mem_238(source_io_mem_238),
    .io_mem_239(source_io_mem_239),
    .io_mem_240(source_io_mem_240),
    .io_mem_241(source_io_mem_241),
    .io_mem_242(source_io_mem_242),
    .io_mem_243(source_io_mem_243),
    .io_mem_244(source_io_mem_244),
    .io_mem_245(source_io_mem_245),
    .io_mem_246(source_io_mem_246),
    .io_mem_247(source_io_mem_247),
    .io_mem_248(source_io_mem_248),
    .io_mem_249(source_io_mem_249),
    .io_mem_250(source_io_mem_250),
    .io_mem_251(source_io_mem_251),
    .io_mem_252(source_io_mem_252),
    .io_mem_253(source_io_mem_253),
    .io_mem_254(source_io_mem_254),
    .io_mem_255(source_io_mem_255),
    .io_sink_reset_n(source_io_sink_reset_n),
    .io_ridx_valid(source_io_ridx_valid),
    .io_widx_valid(source_io_widx_valid)
  );
  AsyncQueueSink sink ( // @[AsyncQueue.scala 156:22]
    .clock(sink_clock),
    .reset(sink_reset),
    .io_deq_ready(sink_io_deq_ready),
    .io_deq_valid(sink_io_deq_valid),
    .io_deq_bits(sink_io_deq_bits),
    .io_ridx(sink_io_ridx),
    .io_widx(sink_io_widx),
    .io_mem_0(sink_io_mem_0),
    .io_mem_1(sink_io_mem_1),
    .io_mem_2(sink_io_mem_2),
    .io_mem_3(sink_io_mem_3),
    .io_mem_4(sink_io_mem_4),
    .io_mem_5(sink_io_mem_5),
    .io_mem_6(sink_io_mem_6),
    .io_mem_7(sink_io_mem_7),
    .io_mem_8(sink_io_mem_8),
    .io_mem_9(sink_io_mem_9),
    .io_mem_10(sink_io_mem_10),
    .io_mem_11(sink_io_mem_11),
    .io_mem_12(sink_io_mem_12),
    .io_mem_13(sink_io_mem_13),
    .io_mem_14(sink_io_mem_14),
    .io_mem_15(sink_io_mem_15),
    .io_mem_16(sink_io_mem_16),
    .io_mem_17(sink_io_mem_17),
    .io_mem_18(sink_io_mem_18),
    .io_mem_19(sink_io_mem_19),
    .io_mem_20(sink_io_mem_20),
    .io_mem_21(sink_io_mem_21),
    .io_mem_22(sink_io_mem_22),
    .io_mem_23(sink_io_mem_23),
    .io_mem_24(sink_io_mem_24),
    .io_mem_25(sink_io_mem_25),
    .io_mem_26(sink_io_mem_26),
    .io_mem_27(sink_io_mem_27),
    .io_mem_28(sink_io_mem_28),
    .io_mem_29(sink_io_mem_29),
    .io_mem_30(sink_io_mem_30),
    .io_mem_31(sink_io_mem_31),
    .io_mem_32(sink_io_mem_32),
    .io_mem_33(sink_io_mem_33),
    .io_mem_34(sink_io_mem_34),
    .io_mem_35(sink_io_mem_35),
    .io_mem_36(sink_io_mem_36),
    .io_mem_37(sink_io_mem_37),
    .io_mem_38(sink_io_mem_38),
    .io_mem_39(sink_io_mem_39),
    .io_mem_40(sink_io_mem_40),
    .io_mem_41(sink_io_mem_41),
    .io_mem_42(sink_io_mem_42),
    .io_mem_43(sink_io_mem_43),
    .io_mem_44(sink_io_mem_44),
    .io_mem_45(sink_io_mem_45),
    .io_mem_46(sink_io_mem_46),
    .io_mem_47(sink_io_mem_47),
    .io_mem_48(sink_io_mem_48),
    .io_mem_49(sink_io_mem_49),
    .io_mem_50(sink_io_mem_50),
    .io_mem_51(sink_io_mem_51),
    .io_mem_52(sink_io_mem_52),
    .io_mem_53(sink_io_mem_53),
    .io_mem_54(sink_io_mem_54),
    .io_mem_55(sink_io_mem_55),
    .io_mem_56(sink_io_mem_56),
    .io_mem_57(sink_io_mem_57),
    .io_mem_58(sink_io_mem_58),
    .io_mem_59(sink_io_mem_59),
    .io_mem_60(sink_io_mem_60),
    .io_mem_61(sink_io_mem_61),
    .io_mem_62(sink_io_mem_62),
    .io_mem_63(sink_io_mem_63),
    .io_mem_64(sink_io_mem_64),
    .io_mem_65(sink_io_mem_65),
    .io_mem_66(sink_io_mem_66),
    .io_mem_67(sink_io_mem_67),
    .io_mem_68(sink_io_mem_68),
    .io_mem_69(sink_io_mem_69),
    .io_mem_70(sink_io_mem_70),
    .io_mem_71(sink_io_mem_71),
    .io_mem_72(sink_io_mem_72),
    .io_mem_73(sink_io_mem_73),
    .io_mem_74(sink_io_mem_74),
    .io_mem_75(sink_io_mem_75),
    .io_mem_76(sink_io_mem_76),
    .io_mem_77(sink_io_mem_77),
    .io_mem_78(sink_io_mem_78),
    .io_mem_79(sink_io_mem_79),
    .io_mem_80(sink_io_mem_80),
    .io_mem_81(sink_io_mem_81),
    .io_mem_82(sink_io_mem_82),
    .io_mem_83(sink_io_mem_83),
    .io_mem_84(sink_io_mem_84),
    .io_mem_85(sink_io_mem_85),
    .io_mem_86(sink_io_mem_86),
    .io_mem_87(sink_io_mem_87),
    .io_mem_88(sink_io_mem_88),
    .io_mem_89(sink_io_mem_89),
    .io_mem_90(sink_io_mem_90),
    .io_mem_91(sink_io_mem_91),
    .io_mem_92(sink_io_mem_92),
    .io_mem_93(sink_io_mem_93),
    .io_mem_94(sink_io_mem_94),
    .io_mem_95(sink_io_mem_95),
    .io_mem_96(sink_io_mem_96),
    .io_mem_97(sink_io_mem_97),
    .io_mem_98(sink_io_mem_98),
    .io_mem_99(sink_io_mem_99),
    .io_mem_100(sink_io_mem_100),
    .io_mem_101(sink_io_mem_101),
    .io_mem_102(sink_io_mem_102),
    .io_mem_103(sink_io_mem_103),
    .io_mem_104(sink_io_mem_104),
    .io_mem_105(sink_io_mem_105),
    .io_mem_106(sink_io_mem_106),
    .io_mem_107(sink_io_mem_107),
    .io_mem_108(sink_io_mem_108),
    .io_mem_109(sink_io_mem_109),
    .io_mem_110(sink_io_mem_110),
    .io_mem_111(sink_io_mem_111),
    .io_mem_112(sink_io_mem_112),
    .io_mem_113(sink_io_mem_113),
    .io_mem_114(sink_io_mem_114),
    .io_mem_115(sink_io_mem_115),
    .io_mem_116(sink_io_mem_116),
    .io_mem_117(sink_io_mem_117),
    .io_mem_118(sink_io_mem_118),
    .io_mem_119(sink_io_mem_119),
    .io_mem_120(sink_io_mem_120),
    .io_mem_121(sink_io_mem_121),
    .io_mem_122(sink_io_mem_122),
    .io_mem_123(sink_io_mem_123),
    .io_mem_124(sink_io_mem_124),
    .io_mem_125(sink_io_mem_125),
    .io_mem_126(sink_io_mem_126),
    .io_mem_127(sink_io_mem_127),
    .io_mem_128(sink_io_mem_128),
    .io_mem_129(sink_io_mem_129),
    .io_mem_130(sink_io_mem_130),
    .io_mem_131(sink_io_mem_131),
    .io_mem_132(sink_io_mem_132),
    .io_mem_133(sink_io_mem_133),
    .io_mem_134(sink_io_mem_134),
    .io_mem_135(sink_io_mem_135),
    .io_mem_136(sink_io_mem_136),
    .io_mem_137(sink_io_mem_137),
    .io_mem_138(sink_io_mem_138),
    .io_mem_139(sink_io_mem_139),
    .io_mem_140(sink_io_mem_140),
    .io_mem_141(sink_io_mem_141),
    .io_mem_142(sink_io_mem_142),
    .io_mem_143(sink_io_mem_143),
    .io_mem_144(sink_io_mem_144),
    .io_mem_145(sink_io_mem_145),
    .io_mem_146(sink_io_mem_146),
    .io_mem_147(sink_io_mem_147),
    .io_mem_148(sink_io_mem_148),
    .io_mem_149(sink_io_mem_149),
    .io_mem_150(sink_io_mem_150),
    .io_mem_151(sink_io_mem_151),
    .io_mem_152(sink_io_mem_152),
    .io_mem_153(sink_io_mem_153),
    .io_mem_154(sink_io_mem_154),
    .io_mem_155(sink_io_mem_155),
    .io_mem_156(sink_io_mem_156),
    .io_mem_157(sink_io_mem_157),
    .io_mem_158(sink_io_mem_158),
    .io_mem_159(sink_io_mem_159),
    .io_mem_160(sink_io_mem_160),
    .io_mem_161(sink_io_mem_161),
    .io_mem_162(sink_io_mem_162),
    .io_mem_163(sink_io_mem_163),
    .io_mem_164(sink_io_mem_164),
    .io_mem_165(sink_io_mem_165),
    .io_mem_166(sink_io_mem_166),
    .io_mem_167(sink_io_mem_167),
    .io_mem_168(sink_io_mem_168),
    .io_mem_169(sink_io_mem_169),
    .io_mem_170(sink_io_mem_170),
    .io_mem_171(sink_io_mem_171),
    .io_mem_172(sink_io_mem_172),
    .io_mem_173(sink_io_mem_173),
    .io_mem_174(sink_io_mem_174),
    .io_mem_175(sink_io_mem_175),
    .io_mem_176(sink_io_mem_176),
    .io_mem_177(sink_io_mem_177),
    .io_mem_178(sink_io_mem_178),
    .io_mem_179(sink_io_mem_179),
    .io_mem_180(sink_io_mem_180),
    .io_mem_181(sink_io_mem_181),
    .io_mem_182(sink_io_mem_182),
    .io_mem_183(sink_io_mem_183),
    .io_mem_184(sink_io_mem_184),
    .io_mem_185(sink_io_mem_185),
    .io_mem_186(sink_io_mem_186),
    .io_mem_187(sink_io_mem_187),
    .io_mem_188(sink_io_mem_188),
    .io_mem_189(sink_io_mem_189),
    .io_mem_190(sink_io_mem_190),
    .io_mem_191(sink_io_mem_191),
    .io_mem_192(sink_io_mem_192),
    .io_mem_193(sink_io_mem_193),
    .io_mem_194(sink_io_mem_194),
    .io_mem_195(sink_io_mem_195),
    .io_mem_196(sink_io_mem_196),
    .io_mem_197(sink_io_mem_197),
    .io_mem_198(sink_io_mem_198),
    .io_mem_199(sink_io_mem_199),
    .io_mem_200(sink_io_mem_200),
    .io_mem_201(sink_io_mem_201),
    .io_mem_202(sink_io_mem_202),
    .io_mem_203(sink_io_mem_203),
    .io_mem_204(sink_io_mem_204),
    .io_mem_205(sink_io_mem_205),
    .io_mem_206(sink_io_mem_206),
    .io_mem_207(sink_io_mem_207),
    .io_mem_208(sink_io_mem_208),
    .io_mem_209(sink_io_mem_209),
    .io_mem_210(sink_io_mem_210),
    .io_mem_211(sink_io_mem_211),
    .io_mem_212(sink_io_mem_212),
    .io_mem_213(sink_io_mem_213),
    .io_mem_214(sink_io_mem_214),
    .io_mem_215(sink_io_mem_215),
    .io_mem_216(sink_io_mem_216),
    .io_mem_217(sink_io_mem_217),
    .io_mem_218(sink_io_mem_218),
    .io_mem_219(sink_io_mem_219),
    .io_mem_220(sink_io_mem_220),
    .io_mem_221(sink_io_mem_221),
    .io_mem_222(sink_io_mem_222),
    .io_mem_223(sink_io_mem_223),
    .io_mem_224(sink_io_mem_224),
    .io_mem_225(sink_io_mem_225),
    .io_mem_226(sink_io_mem_226),
    .io_mem_227(sink_io_mem_227),
    .io_mem_228(sink_io_mem_228),
    .io_mem_229(sink_io_mem_229),
    .io_mem_230(sink_io_mem_230),
    .io_mem_231(sink_io_mem_231),
    .io_mem_232(sink_io_mem_232),
    .io_mem_233(sink_io_mem_233),
    .io_mem_234(sink_io_mem_234),
    .io_mem_235(sink_io_mem_235),
    .io_mem_236(sink_io_mem_236),
    .io_mem_237(sink_io_mem_237),
    .io_mem_238(sink_io_mem_238),
    .io_mem_239(sink_io_mem_239),
    .io_mem_240(sink_io_mem_240),
    .io_mem_241(sink_io_mem_241),
    .io_mem_242(sink_io_mem_242),
    .io_mem_243(sink_io_mem_243),
    .io_mem_244(sink_io_mem_244),
    .io_mem_245(sink_io_mem_245),
    .io_mem_246(sink_io_mem_246),
    .io_mem_247(sink_io_mem_247),
    .io_mem_248(sink_io_mem_248),
    .io_mem_249(sink_io_mem_249),
    .io_mem_250(sink_io_mem_250),
    .io_mem_251(sink_io_mem_251),
    .io_mem_252(sink_io_mem_252),
    .io_mem_253(sink_io_mem_253),
    .io_mem_254(sink_io_mem_254),
    .io_mem_255(sink_io_mem_255),
    .io_source_reset_n(sink_io_source_reset_n),
    .io_ridx_valid(sink_io_ridx_valid),
    .io_widx_valid(sink_io_widx_valid)
  );
  assign io_enq_ready = source_io_enq_ready;
  assign io_deq_valid = sink_io_deq_valid;
  assign io_deq_bits = sink_io_deq_bits;
  assign source_clock = io_enq_clock;
  assign source_reset = 1'h0;
  assign source_io_enq_valid = io_enq_valid;
  assign source_io_enq_bits = io_enq_bits;
  assign source_io_ridx = sink_io_ridx;
  assign source_io_sink_reset_n = 1'h1;
  assign source_io_ridx_valid = sink_io_ridx_valid;
  assign sink_clock = io_deq_clock;
  assign sink_reset = 1'h0;
  assign sink_io_deq_ready = io_deq_ready;
  assign sink_io_widx = source_io_widx;
  assign sink_io_mem_0 = source_io_mem_0;
  assign sink_io_mem_1 = source_io_mem_1;
  assign sink_io_mem_2 = source_io_mem_2;
  assign sink_io_mem_3 = source_io_mem_3;
  assign sink_io_mem_4 = source_io_mem_4;
  assign sink_io_mem_5 = source_io_mem_5;
  assign sink_io_mem_6 = source_io_mem_6;
  assign sink_io_mem_7 = source_io_mem_7;
  assign sink_io_mem_8 = source_io_mem_8;
  assign sink_io_mem_9 = source_io_mem_9;
  assign sink_io_mem_10 = source_io_mem_10;
  assign sink_io_mem_11 = source_io_mem_11;
  assign sink_io_mem_12 = source_io_mem_12;
  assign sink_io_mem_13 = source_io_mem_13;
  assign sink_io_mem_14 = source_io_mem_14;
  assign sink_io_mem_15 = source_io_mem_15;
  assign sink_io_mem_16 = source_io_mem_16;
  assign sink_io_mem_17 = source_io_mem_17;
  assign sink_io_mem_18 = source_io_mem_18;
  assign sink_io_mem_19 = source_io_mem_19;
  assign sink_io_mem_20 = source_io_mem_20;
  assign sink_io_mem_21 = source_io_mem_21;
  assign sink_io_mem_22 = source_io_mem_22;
  assign sink_io_mem_23 = source_io_mem_23;
  assign sink_io_mem_24 = source_io_mem_24;
  assign sink_io_mem_25 = source_io_mem_25;
  assign sink_io_mem_26 = source_io_mem_26;
  assign sink_io_mem_27 = source_io_mem_27;
  assign sink_io_mem_28 = source_io_mem_28;
  assign sink_io_mem_29 = source_io_mem_29;
  assign sink_io_mem_30 = source_io_mem_30;
  assign sink_io_mem_31 = source_io_mem_31;
  assign sink_io_mem_32 = source_io_mem_32;
  assign sink_io_mem_33 = source_io_mem_33;
  assign sink_io_mem_34 = source_io_mem_34;
  assign sink_io_mem_35 = source_io_mem_35;
  assign sink_io_mem_36 = source_io_mem_36;
  assign sink_io_mem_37 = source_io_mem_37;
  assign sink_io_mem_38 = source_io_mem_38;
  assign sink_io_mem_39 = source_io_mem_39;
  assign sink_io_mem_40 = source_io_mem_40;
  assign sink_io_mem_41 = source_io_mem_41;
  assign sink_io_mem_42 = source_io_mem_42;
  assign sink_io_mem_43 = source_io_mem_43;
  assign sink_io_mem_44 = source_io_mem_44;
  assign sink_io_mem_45 = source_io_mem_45;
  assign sink_io_mem_46 = source_io_mem_46;
  assign sink_io_mem_47 = source_io_mem_47;
  assign sink_io_mem_48 = source_io_mem_48;
  assign sink_io_mem_49 = source_io_mem_49;
  assign sink_io_mem_50 = source_io_mem_50;
  assign sink_io_mem_51 = source_io_mem_51;
  assign sink_io_mem_52 = source_io_mem_52;
  assign sink_io_mem_53 = source_io_mem_53;
  assign sink_io_mem_54 = source_io_mem_54;
  assign sink_io_mem_55 = source_io_mem_55;
  assign sink_io_mem_56 = source_io_mem_56;
  assign sink_io_mem_57 = source_io_mem_57;
  assign sink_io_mem_58 = source_io_mem_58;
  assign sink_io_mem_59 = source_io_mem_59;
  assign sink_io_mem_60 = source_io_mem_60;
  assign sink_io_mem_61 = source_io_mem_61;
  assign sink_io_mem_62 = source_io_mem_62;
  assign sink_io_mem_63 = source_io_mem_63;
  assign sink_io_mem_64 = source_io_mem_64;
  assign sink_io_mem_65 = source_io_mem_65;
  assign sink_io_mem_66 = source_io_mem_66;
  assign sink_io_mem_67 = source_io_mem_67;
  assign sink_io_mem_68 = source_io_mem_68;
  assign sink_io_mem_69 = source_io_mem_69;
  assign sink_io_mem_70 = source_io_mem_70;
  assign sink_io_mem_71 = source_io_mem_71;
  assign sink_io_mem_72 = source_io_mem_72;
  assign sink_io_mem_73 = source_io_mem_73;
  assign sink_io_mem_74 = source_io_mem_74;
  assign sink_io_mem_75 = source_io_mem_75;
  assign sink_io_mem_76 = source_io_mem_76;
  assign sink_io_mem_77 = source_io_mem_77;
  assign sink_io_mem_78 = source_io_mem_78;
  assign sink_io_mem_79 = source_io_mem_79;
  assign sink_io_mem_80 = source_io_mem_80;
  assign sink_io_mem_81 = source_io_mem_81;
  assign sink_io_mem_82 = source_io_mem_82;
  assign sink_io_mem_83 = source_io_mem_83;
  assign sink_io_mem_84 = source_io_mem_84;
  assign sink_io_mem_85 = source_io_mem_85;
  assign sink_io_mem_86 = source_io_mem_86;
  assign sink_io_mem_87 = source_io_mem_87;
  assign sink_io_mem_88 = source_io_mem_88;
  assign sink_io_mem_89 = source_io_mem_89;
  assign sink_io_mem_90 = source_io_mem_90;
  assign sink_io_mem_91 = source_io_mem_91;
  assign sink_io_mem_92 = source_io_mem_92;
  assign sink_io_mem_93 = source_io_mem_93;
  assign sink_io_mem_94 = source_io_mem_94;
  assign sink_io_mem_95 = source_io_mem_95;
  assign sink_io_mem_96 = source_io_mem_96;
  assign sink_io_mem_97 = source_io_mem_97;
  assign sink_io_mem_98 = source_io_mem_98;
  assign sink_io_mem_99 = source_io_mem_99;
  assign sink_io_mem_100 = source_io_mem_100;
  assign sink_io_mem_101 = source_io_mem_101;
  assign sink_io_mem_102 = source_io_mem_102;
  assign sink_io_mem_103 = source_io_mem_103;
  assign sink_io_mem_104 = source_io_mem_104;
  assign sink_io_mem_105 = source_io_mem_105;
  assign sink_io_mem_106 = source_io_mem_106;
  assign sink_io_mem_107 = source_io_mem_107;
  assign sink_io_mem_108 = source_io_mem_108;
  assign sink_io_mem_109 = source_io_mem_109;
  assign sink_io_mem_110 = source_io_mem_110;
  assign sink_io_mem_111 = source_io_mem_111;
  assign sink_io_mem_112 = source_io_mem_112;
  assign sink_io_mem_113 = source_io_mem_113;
  assign sink_io_mem_114 = source_io_mem_114;
  assign sink_io_mem_115 = source_io_mem_115;
  assign sink_io_mem_116 = source_io_mem_116;
  assign sink_io_mem_117 = source_io_mem_117;
  assign sink_io_mem_118 = source_io_mem_118;
  assign sink_io_mem_119 = source_io_mem_119;
  assign sink_io_mem_120 = source_io_mem_120;
  assign sink_io_mem_121 = source_io_mem_121;
  assign sink_io_mem_122 = source_io_mem_122;
  assign sink_io_mem_123 = source_io_mem_123;
  assign sink_io_mem_124 = source_io_mem_124;
  assign sink_io_mem_125 = source_io_mem_125;
  assign sink_io_mem_126 = source_io_mem_126;
  assign sink_io_mem_127 = source_io_mem_127;
  assign sink_io_mem_128 = source_io_mem_128;
  assign sink_io_mem_129 = source_io_mem_129;
  assign sink_io_mem_130 = source_io_mem_130;
  assign sink_io_mem_131 = source_io_mem_131;
  assign sink_io_mem_132 = source_io_mem_132;
  assign sink_io_mem_133 = source_io_mem_133;
  assign sink_io_mem_134 = source_io_mem_134;
  assign sink_io_mem_135 = source_io_mem_135;
  assign sink_io_mem_136 = source_io_mem_136;
  assign sink_io_mem_137 = source_io_mem_137;
  assign sink_io_mem_138 = source_io_mem_138;
  assign sink_io_mem_139 = source_io_mem_139;
  assign sink_io_mem_140 = source_io_mem_140;
  assign sink_io_mem_141 = source_io_mem_141;
  assign sink_io_mem_142 = source_io_mem_142;
  assign sink_io_mem_143 = source_io_mem_143;
  assign sink_io_mem_144 = source_io_mem_144;
  assign sink_io_mem_145 = source_io_mem_145;
  assign sink_io_mem_146 = source_io_mem_146;
  assign sink_io_mem_147 = source_io_mem_147;
  assign sink_io_mem_148 = source_io_mem_148;
  assign sink_io_mem_149 = source_io_mem_149;
  assign sink_io_mem_150 = source_io_mem_150;
  assign sink_io_mem_151 = source_io_mem_151;
  assign sink_io_mem_152 = source_io_mem_152;
  assign sink_io_mem_153 = source_io_mem_153;
  assign sink_io_mem_154 = source_io_mem_154;
  assign sink_io_mem_155 = source_io_mem_155;
  assign sink_io_mem_156 = source_io_mem_156;
  assign sink_io_mem_157 = source_io_mem_157;
  assign sink_io_mem_158 = source_io_mem_158;
  assign sink_io_mem_159 = source_io_mem_159;
  assign sink_io_mem_160 = source_io_mem_160;
  assign sink_io_mem_161 = source_io_mem_161;
  assign sink_io_mem_162 = source_io_mem_162;
  assign sink_io_mem_163 = source_io_mem_163;
  assign sink_io_mem_164 = source_io_mem_164;
  assign sink_io_mem_165 = source_io_mem_165;
  assign sink_io_mem_166 = source_io_mem_166;
  assign sink_io_mem_167 = source_io_mem_167;
  assign sink_io_mem_168 = source_io_mem_168;
  assign sink_io_mem_169 = source_io_mem_169;
  assign sink_io_mem_170 = source_io_mem_170;
  assign sink_io_mem_171 = source_io_mem_171;
  assign sink_io_mem_172 = source_io_mem_172;
  assign sink_io_mem_173 = source_io_mem_173;
  assign sink_io_mem_174 = source_io_mem_174;
  assign sink_io_mem_175 = source_io_mem_175;
  assign sink_io_mem_176 = source_io_mem_176;
  assign sink_io_mem_177 = source_io_mem_177;
  assign sink_io_mem_178 = source_io_mem_178;
  assign sink_io_mem_179 = source_io_mem_179;
  assign sink_io_mem_180 = source_io_mem_180;
  assign sink_io_mem_181 = source_io_mem_181;
  assign sink_io_mem_182 = source_io_mem_182;
  assign sink_io_mem_183 = source_io_mem_183;
  assign sink_io_mem_184 = source_io_mem_184;
  assign sink_io_mem_185 = source_io_mem_185;
  assign sink_io_mem_186 = source_io_mem_186;
  assign sink_io_mem_187 = source_io_mem_187;
  assign sink_io_mem_188 = source_io_mem_188;
  assign sink_io_mem_189 = source_io_mem_189;
  assign sink_io_mem_190 = source_io_mem_190;
  assign sink_io_mem_191 = source_io_mem_191;
  assign sink_io_mem_192 = source_io_mem_192;
  assign sink_io_mem_193 = source_io_mem_193;
  assign sink_io_mem_194 = source_io_mem_194;
  assign sink_io_mem_195 = source_io_mem_195;
  assign sink_io_mem_196 = source_io_mem_196;
  assign sink_io_mem_197 = source_io_mem_197;
  assign sink_io_mem_198 = source_io_mem_198;
  assign sink_io_mem_199 = source_io_mem_199;
  assign sink_io_mem_200 = source_io_mem_200;
  assign sink_io_mem_201 = source_io_mem_201;
  assign sink_io_mem_202 = source_io_mem_202;
  assign sink_io_mem_203 = source_io_mem_203;
  assign sink_io_mem_204 = source_io_mem_204;
  assign sink_io_mem_205 = source_io_mem_205;
  assign sink_io_mem_206 = source_io_mem_206;
  assign sink_io_mem_207 = source_io_mem_207;
  assign sink_io_mem_208 = source_io_mem_208;
  assign sink_io_mem_209 = source_io_mem_209;
  assign sink_io_mem_210 = source_io_mem_210;
  assign sink_io_mem_211 = source_io_mem_211;
  assign sink_io_mem_212 = source_io_mem_212;
  assign sink_io_mem_213 = source_io_mem_213;
  assign sink_io_mem_214 = source_io_mem_214;
  assign sink_io_mem_215 = source_io_mem_215;
  assign sink_io_mem_216 = source_io_mem_216;
  assign sink_io_mem_217 = source_io_mem_217;
  assign sink_io_mem_218 = source_io_mem_218;
  assign sink_io_mem_219 = source_io_mem_219;
  assign sink_io_mem_220 = source_io_mem_220;
  assign sink_io_mem_221 = source_io_mem_221;
  assign sink_io_mem_222 = source_io_mem_222;
  assign sink_io_mem_223 = source_io_mem_223;
  assign sink_io_mem_224 = source_io_mem_224;
  assign sink_io_mem_225 = source_io_mem_225;
  assign sink_io_mem_226 = source_io_mem_226;
  assign sink_io_mem_227 = source_io_mem_227;
  assign sink_io_mem_228 = source_io_mem_228;
  assign sink_io_mem_229 = source_io_mem_229;
  assign sink_io_mem_230 = source_io_mem_230;
  assign sink_io_mem_231 = source_io_mem_231;
  assign sink_io_mem_232 = source_io_mem_232;
  assign sink_io_mem_233 = source_io_mem_233;
  assign sink_io_mem_234 = source_io_mem_234;
  assign sink_io_mem_235 = source_io_mem_235;
  assign sink_io_mem_236 = source_io_mem_236;
  assign sink_io_mem_237 = source_io_mem_237;
  assign sink_io_mem_238 = source_io_mem_238;
  assign sink_io_mem_239 = source_io_mem_239;
  assign sink_io_mem_240 = source_io_mem_240;
  assign sink_io_mem_241 = source_io_mem_241;
  assign sink_io_mem_242 = source_io_mem_242;
  assign sink_io_mem_243 = source_io_mem_243;
  assign sink_io_mem_244 = source_io_mem_244;
  assign sink_io_mem_245 = source_io_mem_245;
  assign sink_io_mem_246 = source_io_mem_246;
  assign sink_io_mem_247 = source_io_mem_247;
  assign sink_io_mem_248 = source_io_mem_248;
  assign sink_io_mem_249 = source_io_mem_249;
  assign sink_io_mem_250 = source_io_mem_250;
  assign sink_io_mem_251 = source_io_mem_251;
  assign sink_io_mem_252 = source_io_mem_252;
  assign sink_io_mem_253 = source_io_mem_253;
  assign sink_io_mem_254 = source_io_mem_254;
  assign sink_io_mem_255 = source_io_mem_255;
  assign sink_io_source_reset_n = 1'h1;
  assign sink_io_widx_valid = source_io_widx_valid;
endmodule
module AsyncQueueSource_1(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input  [8:0] io_ridx,
  output [8:0] io_widx,
  output [7:0] io_mem_0,
  output [7:0] io_mem_1,
  output [7:0] io_mem_2,
  output [7:0] io_mem_3,
  output [7:0] io_mem_4,
  output [7:0] io_mem_5,
  output [7:0] io_mem_6,
  output [7:0] io_mem_7,
  output [7:0] io_mem_8,
  output [7:0] io_mem_9,
  output [7:0] io_mem_10,
  output [7:0] io_mem_11,
  output [7:0] io_mem_12,
  output [7:0] io_mem_13,
  output [7:0] io_mem_14,
  output [7:0] io_mem_15,
  output [7:0] io_mem_16,
  output [7:0] io_mem_17,
  output [7:0] io_mem_18,
  output [7:0] io_mem_19,
  output [7:0] io_mem_20,
  output [7:0] io_mem_21,
  output [7:0] io_mem_22,
  output [7:0] io_mem_23,
  output [7:0] io_mem_24,
  output [7:0] io_mem_25,
  output [7:0] io_mem_26,
  output [7:0] io_mem_27,
  output [7:0] io_mem_28,
  output [7:0] io_mem_29,
  output [7:0] io_mem_30,
  output [7:0] io_mem_31,
  output [7:0] io_mem_32,
  output [7:0] io_mem_33,
  output [7:0] io_mem_34,
  output [7:0] io_mem_35,
  output [7:0] io_mem_36,
  output [7:0] io_mem_37,
  output [7:0] io_mem_38,
  output [7:0] io_mem_39,
  output [7:0] io_mem_40,
  output [7:0] io_mem_41,
  output [7:0] io_mem_42,
  output [7:0] io_mem_43,
  output [7:0] io_mem_44,
  output [7:0] io_mem_45,
  output [7:0] io_mem_46,
  output [7:0] io_mem_47,
  output [7:0] io_mem_48,
  output [7:0] io_mem_49,
  output [7:0] io_mem_50,
  output [7:0] io_mem_51,
  output [7:0] io_mem_52,
  output [7:0] io_mem_53,
  output [7:0] io_mem_54,
  output [7:0] io_mem_55,
  output [7:0] io_mem_56,
  output [7:0] io_mem_57,
  output [7:0] io_mem_58,
  output [7:0] io_mem_59,
  output [7:0] io_mem_60,
  output [7:0] io_mem_61,
  output [7:0] io_mem_62,
  output [7:0] io_mem_63,
  output [7:0] io_mem_64,
  output [7:0] io_mem_65,
  output [7:0] io_mem_66,
  output [7:0] io_mem_67,
  output [7:0] io_mem_68,
  output [7:0] io_mem_69,
  output [7:0] io_mem_70,
  output [7:0] io_mem_71,
  output [7:0] io_mem_72,
  output [7:0] io_mem_73,
  output [7:0] io_mem_74,
  output [7:0] io_mem_75,
  output [7:0] io_mem_76,
  output [7:0] io_mem_77,
  output [7:0] io_mem_78,
  output [7:0] io_mem_79,
  output [7:0] io_mem_80,
  output [7:0] io_mem_81,
  output [7:0] io_mem_82,
  output [7:0] io_mem_83,
  output [7:0] io_mem_84,
  output [7:0] io_mem_85,
  output [7:0] io_mem_86,
  output [7:0] io_mem_87,
  output [7:0] io_mem_88,
  output [7:0] io_mem_89,
  output [7:0] io_mem_90,
  output [7:0] io_mem_91,
  output [7:0] io_mem_92,
  output [7:0] io_mem_93,
  output [7:0] io_mem_94,
  output [7:0] io_mem_95,
  output [7:0] io_mem_96,
  output [7:0] io_mem_97,
  output [7:0] io_mem_98,
  output [7:0] io_mem_99,
  output [7:0] io_mem_100,
  output [7:0] io_mem_101,
  output [7:0] io_mem_102,
  output [7:0] io_mem_103,
  output [7:0] io_mem_104,
  output [7:0] io_mem_105,
  output [7:0] io_mem_106,
  output [7:0] io_mem_107,
  output [7:0] io_mem_108,
  output [7:0] io_mem_109,
  output [7:0] io_mem_110,
  output [7:0] io_mem_111,
  output [7:0] io_mem_112,
  output [7:0] io_mem_113,
  output [7:0] io_mem_114,
  output [7:0] io_mem_115,
  output [7:0] io_mem_116,
  output [7:0] io_mem_117,
  output [7:0] io_mem_118,
  output [7:0] io_mem_119,
  output [7:0] io_mem_120,
  output [7:0] io_mem_121,
  output [7:0] io_mem_122,
  output [7:0] io_mem_123,
  output [7:0] io_mem_124,
  output [7:0] io_mem_125,
  output [7:0] io_mem_126,
  output [7:0] io_mem_127,
  output [7:0] io_mem_128,
  output [7:0] io_mem_129,
  output [7:0] io_mem_130,
  output [7:0] io_mem_131,
  output [7:0] io_mem_132,
  output [7:0] io_mem_133,
  output [7:0] io_mem_134,
  output [7:0] io_mem_135,
  output [7:0] io_mem_136,
  output [7:0] io_mem_137,
  output [7:0] io_mem_138,
  output [7:0] io_mem_139,
  output [7:0] io_mem_140,
  output [7:0] io_mem_141,
  output [7:0] io_mem_142,
  output [7:0] io_mem_143,
  output [7:0] io_mem_144,
  output [7:0] io_mem_145,
  output [7:0] io_mem_146,
  output [7:0] io_mem_147,
  output [7:0] io_mem_148,
  output [7:0] io_mem_149,
  output [7:0] io_mem_150,
  output [7:0] io_mem_151,
  output [7:0] io_mem_152,
  output [7:0] io_mem_153,
  output [7:0] io_mem_154,
  output [7:0] io_mem_155,
  output [7:0] io_mem_156,
  output [7:0] io_mem_157,
  output [7:0] io_mem_158,
  output [7:0] io_mem_159,
  output [7:0] io_mem_160,
  output [7:0] io_mem_161,
  output [7:0] io_mem_162,
  output [7:0] io_mem_163,
  output [7:0] io_mem_164,
  output [7:0] io_mem_165,
  output [7:0] io_mem_166,
  output [7:0] io_mem_167,
  output [7:0] io_mem_168,
  output [7:0] io_mem_169,
  output [7:0] io_mem_170,
  output [7:0] io_mem_171,
  output [7:0] io_mem_172,
  output [7:0] io_mem_173,
  output [7:0] io_mem_174,
  output [7:0] io_mem_175,
  output [7:0] io_mem_176,
  output [7:0] io_mem_177,
  output [7:0] io_mem_178,
  output [7:0] io_mem_179,
  output [7:0] io_mem_180,
  output [7:0] io_mem_181,
  output [7:0] io_mem_182,
  output [7:0] io_mem_183,
  output [7:0] io_mem_184,
  output [7:0] io_mem_185,
  output [7:0] io_mem_186,
  output [7:0] io_mem_187,
  output [7:0] io_mem_188,
  output [7:0] io_mem_189,
  output [7:0] io_mem_190,
  output [7:0] io_mem_191,
  output [7:0] io_mem_192,
  output [7:0] io_mem_193,
  output [7:0] io_mem_194,
  output [7:0] io_mem_195,
  output [7:0] io_mem_196,
  output [7:0] io_mem_197,
  output [7:0] io_mem_198,
  output [7:0] io_mem_199,
  output [7:0] io_mem_200,
  output [7:0] io_mem_201,
  output [7:0] io_mem_202,
  output [7:0] io_mem_203,
  output [7:0] io_mem_204,
  output [7:0] io_mem_205,
  output [7:0] io_mem_206,
  output [7:0] io_mem_207,
  output [7:0] io_mem_208,
  output [7:0] io_mem_209,
  output [7:0] io_mem_210,
  output [7:0] io_mem_211,
  output [7:0] io_mem_212,
  output [7:0] io_mem_213,
  output [7:0] io_mem_214,
  output [7:0] io_mem_215,
  output [7:0] io_mem_216,
  output [7:0] io_mem_217,
  output [7:0] io_mem_218,
  output [7:0] io_mem_219,
  output [7:0] io_mem_220,
  output [7:0] io_mem_221,
  output [7:0] io_mem_222,
  output [7:0] io_mem_223,
  output [7:0] io_mem_224,
  output [7:0] io_mem_225,
  output [7:0] io_mem_226,
  output [7:0] io_mem_227,
  output [7:0] io_mem_228,
  output [7:0] io_mem_229,
  output [7:0] io_mem_230,
  output [7:0] io_mem_231,
  output [7:0] io_mem_232,
  output [7:0] io_mem_233,
  output [7:0] io_mem_234,
  output [7:0] io_mem_235,
  output [7:0] io_mem_236,
  output [7:0] io_mem_237,
  output [7:0] io_mem_238,
  output [7:0] io_mem_239,
  output [7:0] io_mem_240,
  output [7:0] io_mem_241,
  output [7:0] io_mem_242,
  output [7:0] io_mem_243,
  output [7:0] io_mem_244,
  output [7:0] io_mem_245,
  output [7:0] io_mem_246,
  output [7:0] io_mem_247,
  output [7:0] io_mem_248,
  output [7:0] io_mem_249,
  output [7:0] io_mem_250,
  output [7:0] io_mem_251,
  output [7:0] io_mem_252,
  output [7:0] io_mem_253,
  output [7:0] io_mem_254,
  output [7:0] io_mem_255,
  input        io_sink_reset_n,
  input        io_ridx_valid,
  output       io_widx_valid
);
  reg [7:0] mem_0; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_0;
  reg [7:0] mem_1; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_1;
  reg [7:0] mem_2; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_2;
  reg [7:0] mem_3; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_3;
  reg [7:0] mem_4; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_4;
  reg [7:0] mem_5; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_5;
  reg [7:0] mem_6; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_6;
  reg [7:0] mem_7; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_7;
  reg [7:0] mem_8; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_8;
  reg [7:0] mem_9; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_9;
  reg [7:0] mem_10; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_10;
  reg [7:0] mem_11; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_11;
  reg [7:0] mem_12; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_12;
  reg [7:0] mem_13; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_13;
  reg [7:0] mem_14; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_14;
  reg [7:0] mem_15; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_15;
  reg [7:0] mem_16; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_16;
  reg [7:0] mem_17; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_17;
  reg [7:0] mem_18; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_18;
  reg [7:0] mem_19; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_19;
  reg [7:0] mem_20; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_20;
  reg [7:0] mem_21; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_21;
  reg [7:0] mem_22; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_22;
  reg [7:0] mem_23; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_23;
  reg [7:0] mem_24; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_24;
  reg [7:0] mem_25; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_25;
  reg [7:0] mem_26; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_26;
  reg [7:0] mem_27; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_27;
  reg [7:0] mem_28; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_28;
  reg [7:0] mem_29; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_29;
  reg [7:0] mem_30; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_30;
  reg [7:0] mem_31; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_31;
  reg [7:0] mem_32; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_32;
  reg [7:0] mem_33; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_33;
  reg [7:0] mem_34; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_34;
  reg [7:0] mem_35; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_35;
  reg [7:0] mem_36; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_36;
  reg [7:0] mem_37; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_37;
  reg [7:0] mem_38; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_38;
  reg [7:0] mem_39; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_39;
  reg [7:0] mem_40; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_40;
  reg [7:0] mem_41; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_41;
  reg [7:0] mem_42; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_42;
  reg [7:0] mem_43; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_43;
  reg [7:0] mem_44; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_44;
  reg [7:0] mem_45; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_45;
  reg [7:0] mem_46; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_46;
  reg [7:0] mem_47; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_47;
  reg [7:0] mem_48; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_48;
  reg [7:0] mem_49; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_49;
  reg [7:0] mem_50; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_50;
  reg [7:0] mem_51; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_51;
  reg [7:0] mem_52; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_52;
  reg [7:0] mem_53; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_53;
  reg [7:0] mem_54; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_54;
  reg [7:0] mem_55; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_55;
  reg [7:0] mem_56; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_56;
  reg [7:0] mem_57; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_57;
  reg [7:0] mem_58; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_58;
  reg [7:0] mem_59; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_59;
  reg [7:0] mem_60; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_60;
  reg [7:0] mem_61; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_61;
  reg [7:0] mem_62; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_62;
  reg [7:0] mem_63; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_63;
  reg [7:0] mem_64; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_64;
  reg [7:0] mem_65; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_65;
  reg [7:0] mem_66; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_66;
  reg [7:0] mem_67; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_67;
  reg [7:0] mem_68; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_68;
  reg [7:0] mem_69; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_69;
  reg [7:0] mem_70; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_70;
  reg [7:0] mem_71; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_71;
  reg [7:0] mem_72; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_72;
  reg [7:0] mem_73; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_73;
  reg [7:0] mem_74; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_74;
  reg [7:0] mem_75; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_75;
  reg [7:0] mem_76; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_76;
  reg [7:0] mem_77; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_77;
  reg [7:0] mem_78; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_78;
  reg [7:0] mem_79; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_79;
  reg [7:0] mem_80; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_80;
  reg [7:0] mem_81; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_81;
  reg [7:0] mem_82; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_82;
  reg [7:0] mem_83; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_83;
  reg [7:0] mem_84; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_84;
  reg [7:0] mem_85; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_85;
  reg [7:0] mem_86; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_86;
  reg [7:0] mem_87; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_87;
  reg [7:0] mem_88; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_88;
  reg [7:0] mem_89; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_89;
  reg [7:0] mem_90; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_90;
  reg [7:0] mem_91; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_91;
  reg [7:0] mem_92; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_92;
  reg [7:0] mem_93; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_93;
  reg [7:0] mem_94; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_94;
  reg [7:0] mem_95; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_95;
  reg [7:0] mem_96; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_96;
  reg [7:0] mem_97; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_97;
  reg [7:0] mem_98; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_98;
  reg [7:0] mem_99; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_99;
  reg [7:0] mem_100; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_100;
  reg [7:0] mem_101; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_101;
  reg [7:0] mem_102; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_102;
  reg [7:0] mem_103; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_103;
  reg [7:0] mem_104; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_104;
  reg [7:0] mem_105; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_105;
  reg [7:0] mem_106; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_106;
  reg [7:0] mem_107; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_107;
  reg [7:0] mem_108; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_108;
  reg [7:0] mem_109; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_109;
  reg [7:0] mem_110; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_110;
  reg [7:0] mem_111; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_111;
  reg [7:0] mem_112; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_112;
  reg [7:0] mem_113; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_113;
  reg [7:0] mem_114; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_114;
  reg [7:0] mem_115; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_115;
  reg [7:0] mem_116; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_116;
  reg [7:0] mem_117; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_117;
  reg [7:0] mem_118; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_118;
  reg [7:0] mem_119; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_119;
  reg [7:0] mem_120; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_120;
  reg [7:0] mem_121; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_121;
  reg [7:0] mem_122; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_122;
  reg [7:0] mem_123; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_123;
  reg [7:0] mem_124; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_124;
  reg [7:0] mem_125; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_125;
  reg [7:0] mem_126; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_126;
  reg [7:0] mem_127; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_127;
  reg [7:0] mem_128; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_128;
  reg [7:0] mem_129; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_129;
  reg [7:0] mem_130; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_130;
  reg [7:0] mem_131; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_131;
  reg [7:0] mem_132; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_132;
  reg [7:0] mem_133; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_133;
  reg [7:0] mem_134; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_134;
  reg [7:0] mem_135; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_135;
  reg [7:0] mem_136; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_136;
  reg [7:0] mem_137; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_137;
  reg [7:0] mem_138; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_138;
  reg [7:0] mem_139; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_139;
  reg [7:0] mem_140; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_140;
  reg [7:0] mem_141; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_141;
  reg [7:0] mem_142; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_142;
  reg [7:0] mem_143; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_143;
  reg [7:0] mem_144; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_144;
  reg [7:0] mem_145; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_145;
  reg [7:0] mem_146; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_146;
  reg [7:0] mem_147; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_147;
  reg [7:0] mem_148; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_148;
  reg [7:0] mem_149; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_149;
  reg [7:0] mem_150; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_150;
  reg [7:0] mem_151; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_151;
  reg [7:0] mem_152; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_152;
  reg [7:0] mem_153; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_153;
  reg [7:0] mem_154; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_154;
  reg [7:0] mem_155; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_155;
  reg [7:0] mem_156; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_156;
  reg [7:0] mem_157; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_157;
  reg [7:0] mem_158; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_158;
  reg [7:0] mem_159; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_159;
  reg [7:0] mem_160; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_160;
  reg [7:0] mem_161; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_161;
  reg [7:0] mem_162; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_162;
  reg [7:0] mem_163; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_163;
  reg [7:0] mem_164; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_164;
  reg [7:0] mem_165; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_165;
  reg [7:0] mem_166; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_166;
  reg [7:0] mem_167; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_167;
  reg [7:0] mem_168; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_168;
  reg [7:0] mem_169; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_169;
  reg [7:0] mem_170; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_170;
  reg [7:0] mem_171; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_171;
  reg [7:0] mem_172; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_172;
  reg [7:0] mem_173; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_173;
  reg [7:0] mem_174; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_174;
  reg [7:0] mem_175; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_175;
  reg [7:0] mem_176; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_176;
  reg [7:0] mem_177; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_177;
  reg [7:0] mem_178; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_178;
  reg [7:0] mem_179; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_179;
  reg [7:0] mem_180; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_180;
  reg [7:0] mem_181; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_181;
  reg [7:0] mem_182; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_182;
  reg [7:0] mem_183; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_183;
  reg [7:0] mem_184; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_184;
  reg [7:0] mem_185; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_185;
  reg [7:0] mem_186; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_186;
  reg [7:0] mem_187; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_187;
  reg [7:0] mem_188; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_188;
  reg [7:0] mem_189; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_189;
  reg [7:0] mem_190; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_190;
  reg [7:0] mem_191; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_191;
  reg [7:0] mem_192; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_192;
  reg [7:0] mem_193; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_193;
  reg [7:0] mem_194; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_194;
  reg [7:0] mem_195; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_195;
  reg [7:0] mem_196; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_196;
  reg [7:0] mem_197; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_197;
  reg [7:0] mem_198; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_198;
  reg [7:0] mem_199; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_199;
  reg [7:0] mem_200; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_200;
  reg [7:0] mem_201; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_201;
  reg [7:0] mem_202; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_202;
  reg [7:0] mem_203; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_203;
  reg [7:0] mem_204; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_204;
  reg [7:0] mem_205; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_205;
  reg [7:0] mem_206; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_206;
  reg [7:0] mem_207; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_207;
  reg [7:0] mem_208; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_208;
  reg [7:0] mem_209; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_209;
  reg [7:0] mem_210; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_210;
  reg [7:0] mem_211; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_211;
  reg [7:0] mem_212; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_212;
  reg [7:0] mem_213; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_213;
  reg [7:0] mem_214; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_214;
  reg [7:0] mem_215; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_215;
  reg [7:0] mem_216; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_216;
  reg [7:0] mem_217; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_217;
  reg [7:0] mem_218; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_218;
  reg [7:0] mem_219; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_219;
  reg [7:0] mem_220; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_220;
  reg [7:0] mem_221; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_221;
  reg [7:0] mem_222; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_222;
  reg [7:0] mem_223; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_223;
  reg [7:0] mem_224; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_224;
  reg [7:0] mem_225; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_225;
  reg [7:0] mem_226; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_226;
  reg [7:0] mem_227; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_227;
  reg [7:0] mem_228; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_228;
  reg [7:0] mem_229; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_229;
  reg [7:0] mem_230; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_230;
  reg [7:0] mem_231; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_231;
  reg [7:0] mem_232; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_232;
  reg [7:0] mem_233; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_233;
  reg [7:0] mem_234; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_234;
  reg [7:0] mem_235; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_235;
  reg [7:0] mem_236; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_236;
  reg [7:0] mem_237; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_237;
  reg [7:0] mem_238; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_238;
  reg [7:0] mem_239; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_239;
  reg [7:0] mem_240; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_240;
  reg [7:0] mem_241; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_241;
  reg [7:0] mem_242; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_242;
  reg [7:0] mem_243; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_243;
  reg [7:0] mem_244; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_244;
  reg [7:0] mem_245; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_245;
  reg [7:0] mem_246; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_246;
  reg [7:0] mem_247; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_247;
  reg [7:0] mem_248; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_248;
  reg [7:0] mem_249; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_249;
  reg [7:0] mem_250; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_250;
  reg [7:0] mem_251; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_251;
  reg [7:0] mem_252; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_252;
  reg [7:0] mem_253; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_253;
  reg [7:0] mem_254; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_254;
  reg [7:0] mem_255; // @[AsyncQueue.scala 41:16]
  reg [31:0] _RAND_255;
  wire  widx_bin_clock; // @[AsyncResetReg.scala 110:21]
  wire  widx_bin_reset; // @[AsyncResetReg.scala 110:21]
  wire [8:0] widx_bin_io_d; // @[AsyncResetReg.scala 110:21]
  wire [8:0] widx_bin_io_q; // @[AsyncResetReg.scala 110:21]
  wire  widx_bin_io_en; // @[AsyncResetReg.scala 110:21]
  wire  ridx_gray_clock; // @[ShiftReg.scala 47:23]
  wire  ridx_gray_reset; // @[ShiftReg.scala 47:23]
  wire [8:0] ridx_gray_io_d; // @[ShiftReg.scala 47:23]
  wire [8:0] ridx_gray_io_q; // @[ShiftReg.scala 47:23]
  wire  ready_reg_clock; // @[AsyncResetReg.scala 110:21]
  wire  ready_reg_reset; // @[AsyncResetReg.scala 110:21]
  wire  ready_reg_io_d; // @[AsyncResetReg.scala 110:21]
  wire  ready_reg_io_q; // @[AsyncResetReg.scala 110:21]
  wire  ready_reg_io_en; // @[AsyncResetReg.scala 110:21]
  wire  widx_gray_clock; // @[AsyncResetReg.scala 110:21]
  wire  widx_gray_reset; // @[AsyncResetReg.scala 110:21]
  wire [8:0] widx_gray_io_d; // @[AsyncResetReg.scala 110:21]
  wire [8:0] widx_gray_io_q; // @[AsyncResetReg.scala 110:21]
  wire  widx_gray_io_en; // @[AsyncResetReg.scala 110:21]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 59:30]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 59:30]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 59:30]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 60:30]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 60:30]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 60:30]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 60:30]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 61:30]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 61:30]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 61:30]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 61:30]
  wire  _T_536; // @[Decoupled.scala 30:37]
  wire  sink_ready;
  wire  _T_538; // @[AsyncQueue.scala 42:49]
  wire [8:0] _GEN_513; // @[AsyncQueue.scala 11:47]
  wire [9:0] _T_543; // @[AsyncQueue.scala 11:47]
  wire [8:0] _T_544; // @[AsyncQueue.scala 11:47]
  wire [8:0] _T_545; // @[AsyncQueue.scala 11:23]
  wire [8:0] _T_547; // @[AsyncQueue.scala 12:32]
  wire [8:0] widx; // @[AsyncQueue.scala 12:17]
  wire [8:0] ridx; // @[ShiftReg.scala 50:24]
  wire [8:0] _T_550; // @[AsyncQueue.scala 44:44]
  wire  _T_551; // @[AsyncQueue.scala 44:34]
  wire  ready; // @[AsyncQueue.scala 44:26]
  wire [7:0] _T_552; // @[AsyncQueue.scala 46:51]
  wire  _T_553; // @[AsyncQueue.scala 46:73]
  wire [7:0] _GEN_514; // @[AsyncQueue.scala 46:86]
  wire [7:0] _T_554; // @[AsyncQueue.scala 46:86]
  wire [7:0] index; // @[AsyncQueue.scala 46:63]
  wire [7:0] _GEN_1; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_2; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_3; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_4; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_5; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_6; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_7; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_8; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_9; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_10; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_11; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_12; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_13; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_14; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_15; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_16; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_17; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_18; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_19; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_20; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_21; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_22; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_23; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_24; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_25; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_26; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_27; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_28; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_29; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_30; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_31; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_32; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_33; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_34; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_35; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_36; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_37; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_38; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_39; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_40; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_41; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_42; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_43; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_44; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_45; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_46; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_47; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_48; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_49; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_50; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_51; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_52; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_53; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_54; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_55; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_56; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_57; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_58; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_59; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_60; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_61; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_62; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_63; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_64; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_65; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_66; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_67; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_68; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_69; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_70; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_71; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_72; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_73; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_74; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_75; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_76; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_77; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_78; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_79; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_80; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_81; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_82; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_83; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_84; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_85; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_86; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_87; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_88; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_89; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_90; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_91; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_92; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_93; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_94; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_95; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_96; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_97; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_98; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_99; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_100; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_101; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_102; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_103; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_104; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_105; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_106; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_107; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_108; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_109; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_110; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_111; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_112; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_113; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_114; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_115; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_116; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_117; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_118; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_119; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_120; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_121; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_122; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_123; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_124; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_125; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_126; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_127; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_128; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_129; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_130; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_131; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_132; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_133; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_134; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_135; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_136; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_137; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_138; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_139; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_140; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_141; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_142; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_143; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_144; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_145; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_146; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_147; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_148; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_149; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_150; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_151; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_152; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_153; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_154; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_155; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_156; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_157; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_158; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_159; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_160; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_161; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_162; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_163; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_164; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_165; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_166; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_167; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_168; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_169; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_170; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_171; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_172; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_173; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_174; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_175; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_176; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_177; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_178; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_179; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_180; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_181; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_182; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_183; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_184; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_185; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_186; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_187; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_188; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_189; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_190; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_191; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_192; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_193; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_194; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_195; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_196; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_197; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_198; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_199; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_200; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_201; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_202; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_203; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_204; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_205; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_206; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_207; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_208; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_209; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_210; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_211; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_212; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_213; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_214; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_215; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_216; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_217; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_218; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_219; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_220; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_221; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_222; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_223; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_224; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_225; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_226; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_227; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_228; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_229; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_230; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_231; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_232; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_233; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_234; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_235; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_236; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_237; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_238; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_239; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_240; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_241; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_242; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_243; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_244; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_245; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_246; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_247; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_248; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_249; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_250; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_251; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_252; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_253; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_254; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_255; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_256; // @[AsyncQueue.scala 47:37]
  wire [7:0] _GEN_257; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_258; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_259; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_260; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_261; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_262; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_263; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_264; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_265; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_266; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_267; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_268; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_269; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_270; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_271; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_272; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_273; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_274; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_275; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_276; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_277; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_278; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_279; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_280; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_281; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_282; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_283; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_284; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_285; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_286; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_287; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_288; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_289; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_290; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_291; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_292; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_293; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_294; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_295; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_296; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_297; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_298; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_299; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_300; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_301; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_302; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_303; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_304; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_305; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_306; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_307; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_308; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_309; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_310; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_311; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_312; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_313; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_314; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_315; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_316; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_317; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_318; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_319; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_320; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_321; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_322; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_323; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_324; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_325; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_326; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_327; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_328; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_329; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_330; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_331; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_332; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_333; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_334; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_335; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_336; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_337; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_338; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_339; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_340; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_341; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_342; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_343; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_344; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_345; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_346; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_347; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_348; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_349; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_350; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_351; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_352; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_353; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_354; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_355; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_356; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_357; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_358; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_359; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_360; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_361; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_362; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_363; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_364; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_365; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_366; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_367; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_368; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_369; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_370; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_371; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_372; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_373; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_374; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_375; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_376; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_377; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_378; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_379; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_380; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_381; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_382; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_383; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_384; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_385; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_386; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_387; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_388; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_389; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_390; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_391; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_392; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_393; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_394; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_395; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_396; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_397; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_398; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_399; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_400; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_401; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_402; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_403; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_404; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_405; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_406; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_407; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_408; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_409; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_410; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_411; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_412; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_413; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_414; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_415; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_416; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_417; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_418; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_419; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_420; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_421; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_422; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_423; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_424; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_425; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_426; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_427; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_428; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_429; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_430; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_431; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_432; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_433; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_434; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_435; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_436; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_437; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_438; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_439; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_440; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_441; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_442; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_443; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_444; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_445; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_446; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_447; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_448; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_449; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_450; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_451; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_452; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_453; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_454; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_455; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_456; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_457; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_458; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_459; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_460; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_461; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_462; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_463; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_464; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_465; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_466; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_467; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_468; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_469; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_470; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_471; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_472; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_473; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_474; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_475; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_476; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_477; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_478; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_479; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_480; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_481; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_482; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_483; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_484; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_485; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_486; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_487; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_488; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_489; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_490; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_491; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_492; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_493; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_494; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_495; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_496; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_497; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_498; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_499; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_500; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_501; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_502; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_503; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_504; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_505; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_506; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_507; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_508; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_509; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_510; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_511; // @[AsyncQueue.scala 47:24]
  wire [7:0] _GEN_512; // @[AsyncQueue.scala 47:24]
  wire  ready_reg_1; // @[AsyncQueue.scala 49:59]
  wire  _T_558; // @[AsyncQueue.scala 50:29]
  wire  _T_563; // @[AsyncQueue.scala 62:36]
  wire  _T_564; // @[AsyncQueue.scala 62:33]
  AsyncResetRegVec_w9_i0 widx_bin ( // @[AsyncResetReg.scala 110:21]
    .clock(widx_bin_clock),
    .reset(widx_bin_reset),
    .io_d(widx_bin_io_d),
    .io_q(widx_bin_io_q),
    .io_en(widx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w9_d3_i0 ridx_gray ( // @[ShiftReg.scala 47:23]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q)
  );
  AsyncResetRegVec_w1_i0 ready_reg ( // @[AsyncResetReg.scala 110:21]
    .clock(ready_reg_clock),
    .reset(ready_reg_reset),
    .io_d(ready_reg_io_d),
    .io_q(ready_reg_io_q),
    .io_en(ready_reg_io_en)
  );
  AsyncResetRegVec_w9_i0 widx_gray ( // @[AsyncResetReg.scala 110:21]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q),
    .io_en(widx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 59:30]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 ( // @[AsyncQueue.scala 60:30]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 ( // @[AsyncQueue.scala 61:30]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  assign _T_536 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 30:37]
  assign sink_ready = AsyncValidSync_2_io_out;
  assign _T_538 = sink_ready == 1'h0; // @[AsyncQueue.scala 42:49]
  assign _GEN_513 = {{8'd0}, _T_536}; // @[AsyncQueue.scala 11:47]
  assign _T_543 = widx_bin_io_q + _GEN_513; // @[AsyncQueue.scala 11:47]
  assign _T_544 = _T_543[8:0]; // @[AsyncQueue.scala 11:47]
  assign _T_545 = _T_538 ? 9'h0 : _T_544; // @[AsyncQueue.scala 11:23]
  assign _T_547 = _T_545 >> 1'h1; // @[AsyncQueue.scala 12:32]
  assign widx = _T_545 ^ _T_547; // @[AsyncQueue.scala 12:17]
  assign ridx = ridx_gray_io_q; // @[ShiftReg.scala 50:24]
  assign _T_550 = ridx ^ 9'h180; // @[AsyncQueue.scala 44:44]
  assign _T_551 = widx != _T_550; // @[AsyncQueue.scala 44:34]
  assign ready = sink_ready & _T_551; // @[AsyncQueue.scala 44:26]
  assign _T_552 = io_widx[7:0]; // @[AsyncQueue.scala 46:51]
  assign _T_553 = io_widx[8]; // @[AsyncQueue.scala 46:73]
  assign _GEN_514 = {{7'd0}, _T_553}; // @[AsyncQueue.scala 46:86]
  assign _T_554 = _GEN_514 << 7; // @[AsyncQueue.scala 46:86]
  assign index = _T_552 ^ _T_554; // @[AsyncQueue.scala 46:63]
  assign _GEN_1 = 8'h0 == index ? io_enq_bits : mem_0; // @[AsyncQueue.scala 47:37]
  assign _GEN_2 = 8'h1 == index ? io_enq_bits : mem_1; // @[AsyncQueue.scala 47:37]
  assign _GEN_3 = 8'h2 == index ? io_enq_bits : mem_2; // @[AsyncQueue.scala 47:37]
  assign _GEN_4 = 8'h3 == index ? io_enq_bits : mem_3; // @[AsyncQueue.scala 47:37]
  assign _GEN_5 = 8'h4 == index ? io_enq_bits : mem_4; // @[AsyncQueue.scala 47:37]
  assign _GEN_6 = 8'h5 == index ? io_enq_bits : mem_5; // @[AsyncQueue.scala 47:37]
  assign _GEN_7 = 8'h6 == index ? io_enq_bits : mem_6; // @[AsyncQueue.scala 47:37]
  assign _GEN_8 = 8'h7 == index ? io_enq_bits : mem_7; // @[AsyncQueue.scala 47:37]
  assign _GEN_9 = 8'h8 == index ? io_enq_bits : mem_8; // @[AsyncQueue.scala 47:37]
  assign _GEN_10 = 8'h9 == index ? io_enq_bits : mem_9; // @[AsyncQueue.scala 47:37]
  assign _GEN_11 = 8'ha == index ? io_enq_bits : mem_10; // @[AsyncQueue.scala 47:37]
  assign _GEN_12 = 8'hb == index ? io_enq_bits : mem_11; // @[AsyncQueue.scala 47:37]
  assign _GEN_13 = 8'hc == index ? io_enq_bits : mem_12; // @[AsyncQueue.scala 47:37]
  assign _GEN_14 = 8'hd == index ? io_enq_bits : mem_13; // @[AsyncQueue.scala 47:37]
  assign _GEN_15 = 8'he == index ? io_enq_bits : mem_14; // @[AsyncQueue.scala 47:37]
  assign _GEN_16 = 8'hf == index ? io_enq_bits : mem_15; // @[AsyncQueue.scala 47:37]
  assign _GEN_17 = 8'h10 == index ? io_enq_bits : mem_16; // @[AsyncQueue.scala 47:37]
  assign _GEN_18 = 8'h11 == index ? io_enq_bits : mem_17; // @[AsyncQueue.scala 47:37]
  assign _GEN_19 = 8'h12 == index ? io_enq_bits : mem_18; // @[AsyncQueue.scala 47:37]
  assign _GEN_20 = 8'h13 == index ? io_enq_bits : mem_19; // @[AsyncQueue.scala 47:37]
  assign _GEN_21 = 8'h14 == index ? io_enq_bits : mem_20; // @[AsyncQueue.scala 47:37]
  assign _GEN_22 = 8'h15 == index ? io_enq_bits : mem_21; // @[AsyncQueue.scala 47:37]
  assign _GEN_23 = 8'h16 == index ? io_enq_bits : mem_22; // @[AsyncQueue.scala 47:37]
  assign _GEN_24 = 8'h17 == index ? io_enq_bits : mem_23; // @[AsyncQueue.scala 47:37]
  assign _GEN_25 = 8'h18 == index ? io_enq_bits : mem_24; // @[AsyncQueue.scala 47:37]
  assign _GEN_26 = 8'h19 == index ? io_enq_bits : mem_25; // @[AsyncQueue.scala 47:37]
  assign _GEN_27 = 8'h1a == index ? io_enq_bits : mem_26; // @[AsyncQueue.scala 47:37]
  assign _GEN_28 = 8'h1b == index ? io_enq_bits : mem_27; // @[AsyncQueue.scala 47:37]
  assign _GEN_29 = 8'h1c == index ? io_enq_bits : mem_28; // @[AsyncQueue.scala 47:37]
  assign _GEN_30 = 8'h1d == index ? io_enq_bits : mem_29; // @[AsyncQueue.scala 47:37]
  assign _GEN_31 = 8'h1e == index ? io_enq_bits : mem_30; // @[AsyncQueue.scala 47:37]
  assign _GEN_32 = 8'h1f == index ? io_enq_bits : mem_31; // @[AsyncQueue.scala 47:37]
  assign _GEN_33 = 8'h20 == index ? io_enq_bits : mem_32; // @[AsyncQueue.scala 47:37]
  assign _GEN_34 = 8'h21 == index ? io_enq_bits : mem_33; // @[AsyncQueue.scala 47:37]
  assign _GEN_35 = 8'h22 == index ? io_enq_bits : mem_34; // @[AsyncQueue.scala 47:37]
  assign _GEN_36 = 8'h23 == index ? io_enq_bits : mem_35; // @[AsyncQueue.scala 47:37]
  assign _GEN_37 = 8'h24 == index ? io_enq_bits : mem_36; // @[AsyncQueue.scala 47:37]
  assign _GEN_38 = 8'h25 == index ? io_enq_bits : mem_37; // @[AsyncQueue.scala 47:37]
  assign _GEN_39 = 8'h26 == index ? io_enq_bits : mem_38; // @[AsyncQueue.scala 47:37]
  assign _GEN_40 = 8'h27 == index ? io_enq_bits : mem_39; // @[AsyncQueue.scala 47:37]
  assign _GEN_41 = 8'h28 == index ? io_enq_bits : mem_40; // @[AsyncQueue.scala 47:37]
  assign _GEN_42 = 8'h29 == index ? io_enq_bits : mem_41; // @[AsyncQueue.scala 47:37]
  assign _GEN_43 = 8'h2a == index ? io_enq_bits : mem_42; // @[AsyncQueue.scala 47:37]
  assign _GEN_44 = 8'h2b == index ? io_enq_bits : mem_43; // @[AsyncQueue.scala 47:37]
  assign _GEN_45 = 8'h2c == index ? io_enq_bits : mem_44; // @[AsyncQueue.scala 47:37]
  assign _GEN_46 = 8'h2d == index ? io_enq_bits : mem_45; // @[AsyncQueue.scala 47:37]
  assign _GEN_47 = 8'h2e == index ? io_enq_bits : mem_46; // @[AsyncQueue.scala 47:37]
  assign _GEN_48 = 8'h2f == index ? io_enq_bits : mem_47; // @[AsyncQueue.scala 47:37]
  assign _GEN_49 = 8'h30 == index ? io_enq_bits : mem_48; // @[AsyncQueue.scala 47:37]
  assign _GEN_50 = 8'h31 == index ? io_enq_bits : mem_49; // @[AsyncQueue.scala 47:37]
  assign _GEN_51 = 8'h32 == index ? io_enq_bits : mem_50; // @[AsyncQueue.scala 47:37]
  assign _GEN_52 = 8'h33 == index ? io_enq_bits : mem_51; // @[AsyncQueue.scala 47:37]
  assign _GEN_53 = 8'h34 == index ? io_enq_bits : mem_52; // @[AsyncQueue.scala 47:37]
  assign _GEN_54 = 8'h35 == index ? io_enq_bits : mem_53; // @[AsyncQueue.scala 47:37]
  assign _GEN_55 = 8'h36 == index ? io_enq_bits : mem_54; // @[AsyncQueue.scala 47:37]
  assign _GEN_56 = 8'h37 == index ? io_enq_bits : mem_55; // @[AsyncQueue.scala 47:37]
  assign _GEN_57 = 8'h38 == index ? io_enq_bits : mem_56; // @[AsyncQueue.scala 47:37]
  assign _GEN_58 = 8'h39 == index ? io_enq_bits : mem_57; // @[AsyncQueue.scala 47:37]
  assign _GEN_59 = 8'h3a == index ? io_enq_bits : mem_58; // @[AsyncQueue.scala 47:37]
  assign _GEN_60 = 8'h3b == index ? io_enq_bits : mem_59; // @[AsyncQueue.scala 47:37]
  assign _GEN_61 = 8'h3c == index ? io_enq_bits : mem_60; // @[AsyncQueue.scala 47:37]
  assign _GEN_62 = 8'h3d == index ? io_enq_bits : mem_61; // @[AsyncQueue.scala 47:37]
  assign _GEN_63 = 8'h3e == index ? io_enq_bits : mem_62; // @[AsyncQueue.scala 47:37]
  assign _GEN_64 = 8'h3f == index ? io_enq_bits : mem_63; // @[AsyncQueue.scala 47:37]
  assign _GEN_65 = 8'h40 == index ? io_enq_bits : mem_64; // @[AsyncQueue.scala 47:37]
  assign _GEN_66 = 8'h41 == index ? io_enq_bits : mem_65; // @[AsyncQueue.scala 47:37]
  assign _GEN_67 = 8'h42 == index ? io_enq_bits : mem_66; // @[AsyncQueue.scala 47:37]
  assign _GEN_68 = 8'h43 == index ? io_enq_bits : mem_67; // @[AsyncQueue.scala 47:37]
  assign _GEN_69 = 8'h44 == index ? io_enq_bits : mem_68; // @[AsyncQueue.scala 47:37]
  assign _GEN_70 = 8'h45 == index ? io_enq_bits : mem_69; // @[AsyncQueue.scala 47:37]
  assign _GEN_71 = 8'h46 == index ? io_enq_bits : mem_70; // @[AsyncQueue.scala 47:37]
  assign _GEN_72 = 8'h47 == index ? io_enq_bits : mem_71; // @[AsyncQueue.scala 47:37]
  assign _GEN_73 = 8'h48 == index ? io_enq_bits : mem_72; // @[AsyncQueue.scala 47:37]
  assign _GEN_74 = 8'h49 == index ? io_enq_bits : mem_73; // @[AsyncQueue.scala 47:37]
  assign _GEN_75 = 8'h4a == index ? io_enq_bits : mem_74; // @[AsyncQueue.scala 47:37]
  assign _GEN_76 = 8'h4b == index ? io_enq_bits : mem_75; // @[AsyncQueue.scala 47:37]
  assign _GEN_77 = 8'h4c == index ? io_enq_bits : mem_76; // @[AsyncQueue.scala 47:37]
  assign _GEN_78 = 8'h4d == index ? io_enq_bits : mem_77; // @[AsyncQueue.scala 47:37]
  assign _GEN_79 = 8'h4e == index ? io_enq_bits : mem_78; // @[AsyncQueue.scala 47:37]
  assign _GEN_80 = 8'h4f == index ? io_enq_bits : mem_79; // @[AsyncQueue.scala 47:37]
  assign _GEN_81 = 8'h50 == index ? io_enq_bits : mem_80; // @[AsyncQueue.scala 47:37]
  assign _GEN_82 = 8'h51 == index ? io_enq_bits : mem_81; // @[AsyncQueue.scala 47:37]
  assign _GEN_83 = 8'h52 == index ? io_enq_bits : mem_82; // @[AsyncQueue.scala 47:37]
  assign _GEN_84 = 8'h53 == index ? io_enq_bits : mem_83; // @[AsyncQueue.scala 47:37]
  assign _GEN_85 = 8'h54 == index ? io_enq_bits : mem_84; // @[AsyncQueue.scala 47:37]
  assign _GEN_86 = 8'h55 == index ? io_enq_bits : mem_85; // @[AsyncQueue.scala 47:37]
  assign _GEN_87 = 8'h56 == index ? io_enq_bits : mem_86; // @[AsyncQueue.scala 47:37]
  assign _GEN_88 = 8'h57 == index ? io_enq_bits : mem_87; // @[AsyncQueue.scala 47:37]
  assign _GEN_89 = 8'h58 == index ? io_enq_bits : mem_88; // @[AsyncQueue.scala 47:37]
  assign _GEN_90 = 8'h59 == index ? io_enq_bits : mem_89; // @[AsyncQueue.scala 47:37]
  assign _GEN_91 = 8'h5a == index ? io_enq_bits : mem_90; // @[AsyncQueue.scala 47:37]
  assign _GEN_92 = 8'h5b == index ? io_enq_bits : mem_91; // @[AsyncQueue.scala 47:37]
  assign _GEN_93 = 8'h5c == index ? io_enq_bits : mem_92; // @[AsyncQueue.scala 47:37]
  assign _GEN_94 = 8'h5d == index ? io_enq_bits : mem_93; // @[AsyncQueue.scala 47:37]
  assign _GEN_95 = 8'h5e == index ? io_enq_bits : mem_94; // @[AsyncQueue.scala 47:37]
  assign _GEN_96 = 8'h5f == index ? io_enq_bits : mem_95; // @[AsyncQueue.scala 47:37]
  assign _GEN_97 = 8'h60 == index ? io_enq_bits : mem_96; // @[AsyncQueue.scala 47:37]
  assign _GEN_98 = 8'h61 == index ? io_enq_bits : mem_97; // @[AsyncQueue.scala 47:37]
  assign _GEN_99 = 8'h62 == index ? io_enq_bits : mem_98; // @[AsyncQueue.scala 47:37]
  assign _GEN_100 = 8'h63 == index ? io_enq_bits : mem_99; // @[AsyncQueue.scala 47:37]
  assign _GEN_101 = 8'h64 == index ? io_enq_bits : mem_100; // @[AsyncQueue.scala 47:37]
  assign _GEN_102 = 8'h65 == index ? io_enq_bits : mem_101; // @[AsyncQueue.scala 47:37]
  assign _GEN_103 = 8'h66 == index ? io_enq_bits : mem_102; // @[AsyncQueue.scala 47:37]
  assign _GEN_104 = 8'h67 == index ? io_enq_bits : mem_103; // @[AsyncQueue.scala 47:37]
  assign _GEN_105 = 8'h68 == index ? io_enq_bits : mem_104; // @[AsyncQueue.scala 47:37]
  assign _GEN_106 = 8'h69 == index ? io_enq_bits : mem_105; // @[AsyncQueue.scala 47:37]
  assign _GEN_107 = 8'h6a == index ? io_enq_bits : mem_106; // @[AsyncQueue.scala 47:37]
  assign _GEN_108 = 8'h6b == index ? io_enq_bits : mem_107; // @[AsyncQueue.scala 47:37]
  assign _GEN_109 = 8'h6c == index ? io_enq_bits : mem_108; // @[AsyncQueue.scala 47:37]
  assign _GEN_110 = 8'h6d == index ? io_enq_bits : mem_109; // @[AsyncQueue.scala 47:37]
  assign _GEN_111 = 8'h6e == index ? io_enq_bits : mem_110; // @[AsyncQueue.scala 47:37]
  assign _GEN_112 = 8'h6f == index ? io_enq_bits : mem_111; // @[AsyncQueue.scala 47:37]
  assign _GEN_113 = 8'h70 == index ? io_enq_bits : mem_112; // @[AsyncQueue.scala 47:37]
  assign _GEN_114 = 8'h71 == index ? io_enq_bits : mem_113; // @[AsyncQueue.scala 47:37]
  assign _GEN_115 = 8'h72 == index ? io_enq_bits : mem_114; // @[AsyncQueue.scala 47:37]
  assign _GEN_116 = 8'h73 == index ? io_enq_bits : mem_115; // @[AsyncQueue.scala 47:37]
  assign _GEN_117 = 8'h74 == index ? io_enq_bits : mem_116; // @[AsyncQueue.scala 47:37]
  assign _GEN_118 = 8'h75 == index ? io_enq_bits : mem_117; // @[AsyncQueue.scala 47:37]
  assign _GEN_119 = 8'h76 == index ? io_enq_bits : mem_118; // @[AsyncQueue.scala 47:37]
  assign _GEN_120 = 8'h77 == index ? io_enq_bits : mem_119; // @[AsyncQueue.scala 47:37]
  assign _GEN_121 = 8'h78 == index ? io_enq_bits : mem_120; // @[AsyncQueue.scala 47:37]
  assign _GEN_122 = 8'h79 == index ? io_enq_bits : mem_121; // @[AsyncQueue.scala 47:37]
  assign _GEN_123 = 8'h7a == index ? io_enq_bits : mem_122; // @[AsyncQueue.scala 47:37]
  assign _GEN_124 = 8'h7b == index ? io_enq_bits : mem_123; // @[AsyncQueue.scala 47:37]
  assign _GEN_125 = 8'h7c == index ? io_enq_bits : mem_124; // @[AsyncQueue.scala 47:37]
  assign _GEN_126 = 8'h7d == index ? io_enq_bits : mem_125; // @[AsyncQueue.scala 47:37]
  assign _GEN_127 = 8'h7e == index ? io_enq_bits : mem_126; // @[AsyncQueue.scala 47:37]
  assign _GEN_128 = 8'h7f == index ? io_enq_bits : mem_127; // @[AsyncQueue.scala 47:37]
  assign _GEN_129 = 8'h80 == index ? io_enq_bits : mem_128; // @[AsyncQueue.scala 47:37]
  assign _GEN_130 = 8'h81 == index ? io_enq_bits : mem_129; // @[AsyncQueue.scala 47:37]
  assign _GEN_131 = 8'h82 == index ? io_enq_bits : mem_130; // @[AsyncQueue.scala 47:37]
  assign _GEN_132 = 8'h83 == index ? io_enq_bits : mem_131; // @[AsyncQueue.scala 47:37]
  assign _GEN_133 = 8'h84 == index ? io_enq_bits : mem_132; // @[AsyncQueue.scala 47:37]
  assign _GEN_134 = 8'h85 == index ? io_enq_bits : mem_133; // @[AsyncQueue.scala 47:37]
  assign _GEN_135 = 8'h86 == index ? io_enq_bits : mem_134; // @[AsyncQueue.scala 47:37]
  assign _GEN_136 = 8'h87 == index ? io_enq_bits : mem_135; // @[AsyncQueue.scala 47:37]
  assign _GEN_137 = 8'h88 == index ? io_enq_bits : mem_136; // @[AsyncQueue.scala 47:37]
  assign _GEN_138 = 8'h89 == index ? io_enq_bits : mem_137; // @[AsyncQueue.scala 47:37]
  assign _GEN_139 = 8'h8a == index ? io_enq_bits : mem_138; // @[AsyncQueue.scala 47:37]
  assign _GEN_140 = 8'h8b == index ? io_enq_bits : mem_139; // @[AsyncQueue.scala 47:37]
  assign _GEN_141 = 8'h8c == index ? io_enq_bits : mem_140; // @[AsyncQueue.scala 47:37]
  assign _GEN_142 = 8'h8d == index ? io_enq_bits : mem_141; // @[AsyncQueue.scala 47:37]
  assign _GEN_143 = 8'h8e == index ? io_enq_bits : mem_142; // @[AsyncQueue.scala 47:37]
  assign _GEN_144 = 8'h8f == index ? io_enq_bits : mem_143; // @[AsyncQueue.scala 47:37]
  assign _GEN_145 = 8'h90 == index ? io_enq_bits : mem_144; // @[AsyncQueue.scala 47:37]
  assign _GEN_146 = 8'h91 == index ? io_enq_bits : mem_145; // @[AsyncQueue.scala 47:37]
  assign _GEN_147 = 8'h92 == index ? io_enq_bits : mem_146; // @[AsyncQueue.scala 47:37]
  assign _GEN_148 = 8'h93 == index ? io_enq_bits : mem_147; // @[AsyncQueue.scala 47:37]
  assign _GEN_149 = 8'h94 == index ? io_enq_bits : mem_148; // @[AsyncQueue.scala 47:37]
  assign _GEN_150 = 8'h95 == index ? io_enq_bits : mem_149; // @[AsyncQueue.scala 47:37]
  assign _GEN_151 = 8'h96 == index ? io_enq_bits : mem_150; // @[AsyncQueue.scala 47:37]
  assign _GEN_152 = 8'h97 == index ? io_enq_bits : mem_151; // @[AsyncQueue.scala 47:37]
  assign _GEN_153 = 8'h98 == index ? io_enq_bits : mem_152; // @[AsyncQueue.scala 47:37]
  assign _GEN_154 = 8'h99 == index ? io_enq_bits : mem_153; // @[AsyncQueue.scala 47:37]
  assign _GEN_155 = 8'h9a == index ? io_enq_bits : mem_154; // @[AsyncQueue.scala 47:37]
  assign _GEN_156 = 8'h9b == index ? io_enq_bits : mem_155; // @[AsyncQueue.scala 47:37]
  assign _GEN_157 = 8'h9c == index ? io_enq_bits : mem_156; // @[AsyncQueue.scala 47:37]
  assign _GEN_158 = 8'h9d == index ? io_enq_bits : mem_157; // @[AsyncQueue.scala 47:37]
  assign _GEN_159 = 8'h9e == index ? io_enq_bits : mem_158; // @[AsyncQueue.scala 47:37]
  assign _GEN_160 = 8'h9f == index ? io_enq_bits : mem_159; // @[AsyncQueue.scala 47:37]
  assign _GEN_161 = 8'ha0 == index ? io_enq_bits : mem_160; // @[AsyncQueue.scala 47:37]
  assign _GEN_162 = 8'ha1 == index ? io_enq_bits : mem_161; // @[AsyncQueue.scala 47:37]
  assign _GEN_163 = 8'ha2 == index ? io_enq_bits : mem_162; // @[AsyncQueue.scala 47:37]
  assign _GEN_164 = 8'ha3 == index ? io_enq_bits : mem_163; // @[AsyncQueue.scala 47:37]
  assign _GEN_165 = 8'ha4 == index ? io_enq_bits : mem_164; // @[AsyncQueue.scala 47:37]
  assign _GEN_166 = 8'ha5 == index ? io_enq_bits : mem_165; // @[AsyncQueue.scala 47:37]
  assign _GEN_167 = 8'ha6 == index ? io_enq_bits : mem_166; // @[AsyncQueue.scala 47:37]
  assign _GEN_168 = 8'ha7 == index ? io_enq_bits : mem_167; // @[AsyncQueue.scala 47:37]
  assign _GEN_169 = 8'ha8 == index ? io_enq_bits : mem_168; // @[AsyncQueue.scala 47:37]
  assign _GEN_170 = 8'ha9 == index ? io_enq_bits : mem_169; // @[AsyncQueue.scala 47:37]
  assign _GEN_171 = 8'haa == index ? io_enq_bits : mem_170; // @[AsyncQueue.scala 47:37]
  assign _GEN_172 = 8'hab == index ? io_enq_bits : mem_171; // @[AsyncQueue.scala 47:37]
  assign _GEN_173 = 8'hac == index ? io_enq_bits : mem_172; // @[AsyncQueue.scala 47:37]
  assign _GEN_174 = 8'had == index ? io_enq_bits : mem_173; // @[AsyncQueue.scala 47:37]
  assign _GEN_175 = 8'hae == index ? io_enq_bits : mem_174; // @[AsyncQueue.scala 47:37]
  assign _GEN_176 = 8'haf == index ? io_enq_bits : mem_175; // @[AsyncQueue.scala 47:37]
  assign _GEN_177 = 8'hb0 == index ? io_enq_bits : mem_176; // @[AsyncQueue.scala 47:37]
  assign _GEN_178 = 8'hb1 == index ? io_enq_bits : mem_177; // @[AsyncQueue.scala 47:37]
  assign _GEN_179 = 8'hb2 == index ? io_enq_bits : mem_178; // @[AsyncQueue.scala 47:37]
  assign _GEN_180 = 8'hb3 == index ? io_enq_bits : mem_179; // @[AsyncQueue.scala 47:37]
  assign _GEN_181 = 8'hb4 == index ? io_enq_bits : mem_180; // @[AsyncQueue.scala 47:37]
  assign _GEN_182 = 8'hb5 == index ? io_enq_bits : mem_181; // @[AsyncQueue.scala 47:37]
  assign _GEN_183 = 8'hb6 == index ? io_enq_bits : mem_182; // @[AsyncQueue.scala 47:37]
  assign _GEN_184 = 8'hb7 == index ? io_enq_bits : mem_183; // @[AsyncQueue.scala 47:37]
  assign _GEN_185 = 8'hb8 == index ? io_enq_bits : mem_184; // @[AsyncQueue.scala 47:37]
  assign _GEN_186 = 8'hb9 == index ? io_enq_bits : mem_185; // @[AsyncQueue.scala 47:37]
  assign _GEN_187 = 8'hba == index ? io_enq_bits : mem_186; // @[AsyncQueue.scala 47:37]
  assign _GEN_188 = 8'hbb == index ? io_enq_bits : mem_187; // @[AsyncQueue.scala 47:37]
  assign _GEN_189 = 8'hbc == index ? io_enq_bits : mem_188; // @[AsyncQueue.scala 47:37]
  assign _GEN_190 = 8'hbd == index ? io_enq_bits : mem_189; // @[AsyncQueue.scala 47:37]
  assign _GEN_191 = 8'hbe == index ? io_enq_bits : mem_190; // @[AsyncQueue.scala 47:37]
  assign _GEN_192 = 8'hbf == index ? io_enq_bits : mem_191; // @[AsyncQueue.scala 47:37]
  assign _GEN_193 = 8'hc0 == index ? io_enq_bits : mem_192; // @[AsyncQueue.scala 47:37]
  assign _GEN_194 = 8'hc1 == index ? io_enq_bits : mem_193; // @[AsyncQueue.scala 47:37]
  assign _GEN_195 = 8'hc2 == index ? io_enq_bits : mem_194; // @[AsyncQueue.scala 47:37]
  assign _GEN_196 = 8'hc3 == index ? io_enq_bits : mem_195; // @[AsyncQueue.scala 47:37]
  assign _GEN_197 = 8'hc4 == index ? io_enq_bits : mem_196; // @[AsyncQueue.scala 47:37]
  assign _GEN_198 = 8'hc5 == index ? io_enq_bits : mem_197; // @[AsyncQueue.scala 47:37]
  assign _GEN_199 = 8'hc6 == index ? io_enq_bits : mem_198; // @[AsyncQueue.scala 47:37]
  assign _GEN_200 = 8'hc7 == index ? io_enq_bits : mem_199; // @[AsyncQueue.scala 47:37]
  assign _GEN_201 = 8'hc8 == index ? io_enq_bits : mem_200; // @[AsyncQueue.scala 47:37]
  assign _GEN_202 = 8'hc9 == index ? io_enq_bits : mem_201; // @[AsyncQueue.scala 47:37]
  assign _GEN_203 = 8'hca == index ? io_enq_bits : mem_202; // @[AsyncQueue.scala 47:37]
  assign _GEN_204 = 8'hcb == index ? io_enq_bits : mem_203; // @[AsyncQueue.scala 47:37]
  assign _GEN_205 = 8'hcc == index ? io_enq_bits : mem_204; // @[AsyncQueue.scala 47:37]
  assign _GEN_206 = 8'hcd == index ? io_enq_bits : mem_205; // @[AsyncQueue.scala 47:37]
  assign _GEN_207 = 8'hce == index ? io_enq_bits : mem_206; // @[AsyncQueue.scala 47:37]
  assign _GEN_208 = 8'hcf == index ? io_enq_bits : mem_207; // @[AsyncQueue.scala 47:37]
  assign _GEN_209 = 8'hd0 == index ? io_enq_bits : mem_208; // @[AsyncQueue.scala 47:37]
  assign _GEN_210 = 8'hd1 == index ? io_enq_bits : mem_209; // @[AsyncQueue.scala 47:37]
  assign _GEN_211 = 8'hd2 == index ? io_enq_bits : mem_210; // @[AsyncQueue.scala 47:37]
  assign _GEN_212 = 8'hd3 == index ? io_enq_bits : mem_211; // @[AsyncQueue.scala 47:37]
  assign _GEN_213 = 8'hd4 == index ? io_enq_bits : mem_212; // @[AsyncQueue.scala 47:37]
  assign _GEN_214 = 8'hd5 == index ? io_enq_bits : mem_213; // @[AsyncQueue.scala 47:37]
  assign _GEN_215 = 8'hd6 == index ? io_enq_bits : mem_214; // @[AsyncQueue.scala 47:37]
  assign _GEN_216 = 8'hd7 == index ? io_enq_bits : mem_215; // @[AsyncQueue.scala 47:37]
  assign _GEN_217 = 8'hd8 == index ? io_enq_bits : mem_216; // @[AsyncQueue.scala 47:37]
  assign _GEN_218 = 8'hd9 == index ? io_enq_bits : mem_217; // @[AsyncQueue.scala 47:37]
  assign _GEN_219 = 8'hda == index ? io_enq_bits : mem_218; // @[AsyncQueue.scala 47:37]
  assign _GEN_220 = 8'hdb == index ? io_enq_bits : mem_219; // @[AsyncQueue.scala 47:37]
  assign _GEN_221 = 8'hdc == index ? io_enq_bits : mem_220; // @[AsyncQueue.scala 47:37]
  assign _GEN_222 = 8'hdd == index ? io_enq_bits : mem_221; // @[AsyncQueue.scala 47:37]
  assign _GEN_223 = 8'hde == index ? io_enq_bits : mem_222; // @[AsyncQueue.scala 47:37]
  assign _GEN_224 = 8'hdf == index ? io_enq_bits : mem_223; // @[AsyncQueue.scala 47:37]
  assign _GEN_225 = 8'he0 == index ? io_enq_bits : mem_224; // @[AsyncQueue.scala 47:37]
  assign _GEN_226 = 8'he1 == index ? io_enq_bits : mem_225; // @[AsyncQueue.scala 47:37]
  assign _GEN_227 = 8'he2 == index ? io_enq_bits : mem_226; // @[AsyncQueue.scala 47:37]
  assign _GEN_228 = 8'he3 == index ? io_enq_bits : mem_227; // @[AsyncQueue.scala 47:37]
  assign _GEN_229 = 8'he4 == index ? io_enq_bits : mem_228; // @[AsyncQueue.scala 47:37]
  assign _GEN_230 = 8'he5 == index ? io_enq_bits : mem_229; // @[AsyncQueue.scala 47:37]
  assign _GEN_231 = 8'he6 == index ? io_enq_bits : mem_230; // @[AsyncQueue.scala 47:37]
  assign _GEN_232 = 8'he7 == index ? io_enq_bits : mem_231; // @[AsyncQueue.scala 47:37]
  assign _GEN_233 = 8'he8 == index ? io_enq_bits : mem_232; // @[AsyncQueue.scala 47:37]
  assign _GEN_234 = 8'he9 == index ? io_enq_bits : mem_233; // @[AsyncQueue.scala 47:37]
  assign _GEN_235 = 8'hea == index ? io_enq_bits : mem_234; // @[AsyncQueue.scala 47:37]
  assign _GEN_236 = 8'heb == index ? io_enq_bits : mem_235; // @[AsyncQueue.scala 47:37]
  assign _GEN_237 = 8'hec == index ? io_enq_bits : mem_236; // @[AsyncQueue.scala 47:37]
  assign _GEN_238 = 8'hed == index ? io_enq_bits : mem_237; // @[AsyncQueue.scala 47:37]
  assign _GEN_239 = 8'hee == index ? io_enq_bits : mem_238; // @[AsyncQueue.scala 47:37]
  assign _GEN_240 = 8'hef == index ? io_enq_bits : mem_239; // @[AsyncQueue.scala 47:37]
  assign _GEN_241 = 8'hf0 == index ? io_enq_bits : mem_240; // @[AsyncQueue.scala 47:37]
  assign _GEN_242 = 8'hf1 == index ? io_enq_bits : mem_241; // @[AsyncQueue.scala 47:37]
  assign _GEN_243 = 8'hf2 == index ? io_enq_bits : mem_242; // @[AsyncQueue.scala 47:37]
  assign _GEN_244 = 8'hf3 == index ? io_enq_bits : mem_243; // @[AsyncQueue.scala 47:37]
  assign _GEN_245 = 8'hf4 == index ? io_enq_bits : mem_244; // @[AsyncQueue.scala 47:37]
  assign _GEN_246 = 8'hf5 == index ? io_enq_bits : mem_245; // @[AsyncQueue.scala 47:37]
  assign _GEN_247 = 8'hf6 == index ? io_enq_bits : mem_246; // @[AsyncQueue.scala 47:37]
  assign _GEN_248 = 8'hf7 == index ? io_enq_bits : mem_247; // @[AsyncQueue.scala 47:37]
  assign _GEN_249 = 8'hf8 == index ? io_enq_bits : mem_248; // @[AsyncQueue.scala 47:37]
  assign _GEN_250 = 8'hf9 == index ? io_enq_bits : mem_249; // @[AsyncQueue.scala 47:37]
  assign _GEN_251 = 8'hfa == index ? io_enq_bits : mem_250; // @[AsyncQueue.scala 47:37]
  assign _GEN_252 = 8'hfb == index ? io_enq_bits : mem_251; // @[AsyncQueue.scala 47:37]
  assign _GEN_253 = 8'hfc == index ? io_enq_bits : mem_252; // @[AsyncQueue.scala 47:37]
  assign _GEN_254 = 8'hfd == index ? io_enq_bits : mem_253; // @[AsyncQueue.scala 47:37]
  assign _GEN_255 = 8'hfe == index ? io_enq_bits : mem_254; // @[AsyncQueue.scala 47:37]
  assign _GEN_256 = 8'hff == index ? io_enq_bits : mem_255; // @[AsyncQueue.scala 47:37]
  assign _GEN_257 = _T_536 ? _GEN_1 : mem_0; // @[AsyncQueue.scala 47:24]
  assign _GEN_258 = _T_536 ? _GEN_2 : mem_1; // @[AsyncQueue.scala 47:24]
  assign _GEN_259 = _T_536 ? _GEN_3 : mem_2; // @[AsyncQueue.scala 47:24]
  assign _GEN_260 = _T_536 ? _GEN_4 : mem_3; // @[AsyncQueue.scala 47:24]
  assign _GEN_261 = _T_536 ? _GEN_5 : mem_4; // @[AsyncQueue.scala 47:24]
  assign _GEN_262 = _T_536 ? _GEN_6 : mem_5; // @[AsyncQueue.scala 47:24]
  assign _GEN_263 = _T_536 ? _GEN_7 : mem_6; // @[AsyncQueue.scala 47:24]
  assign _GEN_264 = _T_536 ? _GEN_8 : mem_7; // @[AsyncQueue.scala 47:24]
  assign _GEN_265 = _T_536 ? _GEN_9 : mem_8; // @[AsyncQueue.scala 47:24]
  assign _GEN_266 = _T_536 ? _GEN_10 : mem_9; // @[AsyncQueue.scala 47:24]
  assign _GEN_267 = _T_536 ? _GEN_11 : mem_10; // @[AsyncQueue.scala 47:24]
  assign _GEN_268 = _T_536 ? _GEN_12 : mem_11; // @[AsyncQueue.scala 47:24]
  assign _GEN_269 = _T_536 ? _GEN_13 : mem_12; // @[AsyncQueue.scala 47:24]
  assign _GEN_270 = _T_536 ? _GEN_14 : mem_13; // @[AsyncQueue.scala 47:24]
  assign _GEN_271 = _T_536 ? _GEN_15 : mem_14; // @[AsyncQueue.scala 47:24]
  assign _GEN_272 = _T_536 ? _GEN_16 : mem_15; // @[AsyncQueue.scala 47:24]
  assign _GEN_273 = _T_536 ? _GEN_17 : mem_16; // @[AsyncQueue.scala 47:24]
  assign _GEN_274 = _T_536 ? _GEN_18 : mem_17; // @[AsyncQueue.scala 47:24]
  assign _GEN_275 = _T_536 ? _GEN_19 : mem_18; // @[AsyncQueue.scala 47:24]
  assign _GEN_276 = _T_536 ? _GEN_20 : mem_19; // @[AsyncQueue.scala 47:24]
  assign _GEN_277 = _T_536 ? _GEN_21 : mem_20; // @[AsyncQueue.scala 47:24]
  assign _GEN_278 = _T_536 ? _GEN_22 : mem_21; // @[AsyncQueue.scala 47:24]
  assign _GEN_279 = _T_536 ? _GEN_23 : mem_22; // @[AsyncQueue.scala 47:24]
  assign _GEN_280 = _T_536 ? _GEN_24 : mem_23; // @[AsyncQueue.scala 47:24]
  assign _GEN_281 = _T_536 ? _GEN_25 : mem_24; // @[AsyncQueue.scala 47:24]
  assign _GEN_282 = _T_536 ? _GEN_26 : mem_25; // @[AsyncQueue.scala 47:24]
  assign _GEN_283 = _T_536 ? _GEN_27 : mem_26; // @[AsyncQueue.scala 47:24]
  assign _GEN_284 = _T_536 ? _GEN_28 : mem_27; // @[AsyncQueue.scala 47:24]
  assign _GEN_285 = _T_536 ? _GEN_29 : mem_28; // @[AsyncQueue.scala 47:24]
  assign _GEN_286 = _T_536 ? _GEN_30 : mem_29; // @[AsyncQueue.scala 47:24]
  assign _GEN_287 = _T_536 ? _GEN_31 : mem_30; // @[AsyncQueue.scala 47:24]
  assign _GEN_288 = _T_536 ? _GEN_32 : mem_31; // @[AsyncQueue.scala 47:24]
  assign _GEN_289 = _T_536 ? _GEN_33 : mem_32; // @[AsyncQueue.scala 47:24]
  assign _GEN_290 = _T_536 ? _GEN_34 : mem_33; // @[AsyncQueue.scala 47:24]
  assign _GEN_291 = _T_536 ? _GEN_35 : mem_34; // @[AsyncQueue.scala 47:24]
  assign _GEN_292 = _T_536 ? _GEN_36 : mem_35; // @[AsyncQueue.scala 47:24]
  assign _GEN_293 = _T_536 ? _GEN_37 : mem_36; // @[AsyncQueue.scala 47:24]
  assign _GEN_294 = _T_536 ? _GEN_38 : mem_37; // @[AsyncQueue.scala 47:24]
  assign _GEN_295 = _T_536 ? _GEN_39 : mem_38; // @[AsyncQueue.scala 47:24]
  assign _GEN_296 = _T_536 ? _GEN_40 : mem_39; // @[AsyncQueue.scala 47:24]
  assign _GEN_297 = _T_536 ? _GEN_41 : mem_40; // @[AsyncQueue.scala 47:24]
  assign _GEN_298 = _T_536 ? _GEN_42 : mem_41; // @[AsyncQueue.scala 47:24]
  assign _GEN_299 = _T_536 ? _GEN_43 : mem_42; // @[AsyncQueue.scala 47:24]
  assign _GEN_300 = _T_536 ? _GEN_44 : mem_43; // @[AsyncQueue.scala 47:24]
  assign _GEN_301 = _T_536 ? _GEN_45 : mem_44; // @[AsyncQueue.scala 47:24]
  assign _GEN_302 = _T_536 ? _GEN_46 : mem_45; // @[AsyncQueue.scala 47:24]
  assign _GEN_303 = _T_536 ? _GEN_47 : mem_46; // @[AsyncQueue.scala 47:24]
  assign _GEN_304 = _T_536 ? _GEN_48 : mem_47; // @[AsyncQueue.scala 47:24]
  assign _GEN_305 = _T_536 ? _GEN_49 : mem_48; // @[AsyncQueue.scala 47:24]
  assign _GEN_306 = _T_536 ? _GEN_50 : mem_49; // @[AsyncQueue.scala 47:24]
  assign _GEN_307 = _T_536 ? _GEN_51 : mem_50; // @[AsyncQueue.scala 47:24]
  assign _GEN_308 = _T_536 ? _GEN_52 : mem_51; // @[AsyncQueue.scala 47:24]
  assign _GEN_309 = _T_536 ? _GEN_53 : mem_52; // @[AsyncQueue.scala 47:24]
  assign _GEN_310 = _T_536 ? _GEN_54 : mem_53; // @[AsyncQueue.scala 47:24]
  assign _GEN_311 = _T_536 ? _GEN_55 : mem_54; // @[AsyncQueue.scala 47:24]
  assign _GEN_312 = _T_536 ? _GEN_56 : mem_55; // @[AsyncQueue.scala 47:24]
  assign _GEN_313 = _T_536 ? _GEN_57 : mem_56; // @[AsyncQueue.scala 47:24]
  assign _GEN_314 = _T_536 ? _GEN_58 : mem_57; // @[AsyncQueue.scala 47:24]
  assign _GEN_315 = _T_536 ? _GEN_59 : mem_58; // @[AsyncQueue.scala 47:24]
  assign _GEN_316 = _T_536 ? _GEN_60 : mem_59; // @[AsyncQueue.scala 47:24]
  assign _GEN_317 = _T_536 ? _GEN_61 : mem_60; // @[AsyncQueue.scala 47:24]
  assign _GEN_318 = _T_536 ? _GEN_62 : mem_61; // @[AsyncQueue.scala 47:24]
  assign _GEN_319 = _T_536 ? _GEN_63 : mem_62; // @[AsyncQueue.scala 47:24]
  assign _GEN_320 = _T_536 ? _GEN_64 : mem_63; // @[AsyncQueue.scala 47:24]
  assign _GEN_321 = _T_536 ? _GEN_65 : mem_64; // @[AsyncQueue.scala 47:24]
  assign _GEN_322 = _T_536 ? _GEN_66 : mem_65; // @[AsyncQueue.scala 47:24]
  assign _GEN_323 = _T_536 ? _GEN_67 : mem_66; // @[AsyncQueue.scala 47:24]
  assign _GEN_324 = _T_536 ? _GEN_68 : mem_67; // @[AsyncQueue.scala 47:24]
  assign _GEN_325 = _T_536 ? _GEN_69 : mem_68; // @[AsyncQueue.scala 47:24]
  assign _GEN_326 = _T_536 ? _GEN_70 : mem_69; // @[AsyncQueue.scala 47:24]
  assign _GEN_327 = _T_536 ? _GEN_71 : mem_70; // @[AsyncQueue.scala 47:24]
  assign _GEN_328 = _T_536 ? _GEN_72 : mem_71; // @[AsyncQueue.scala 47:24]
  assign _GEN_329 = _T_536 ? _GEN_73 : mem_72; // @[AsyncQueue.scala 47:24]
  assign _GEN_330 = _T_536 ? _GEN_74 : mem_73; // @[AsyncQueue.scala 47:24]
  assign _GEN_331 = _T_536 ? _GEN_75 : mem_74; // @[AsyncQueue.scala 47:24]
  assign _GEN_332 = _T_536 ? _GEN_76 : mem_75; // @[AsyncQueue.scala 47:24]
  assign _GEN_333 = _T_536 ? _GEN_77 : mem_76; // @[AsyncQueue.scala 47:24]
  assign _GEN_334 = _T_536 ? _GEN_78 : mem_77; // @[AsyncQueue.scala 47:24]
  assign _GEN_335 = _T_536 ? _GEN_79 : mem_78; // @[AsyncQueue.scala 47:24]
  assign _GEN_336 = _T_536 ? _GEN_80 : mem_79; // @[AsyncQueue.scala 47:24]
  assign _GEN_337 = _T_536 ? _GEN_81 : mem_80; // @[AsyncQueue.scala 47:24]
  assign _GEN_338 = _T_536 ? _GEN_82 : mem_81; // @[AsyncQueue.scala 47:24]
  assign _GEN_339 = _T_536 ? _GEN_83 : mem_82; // @[AsyncQueue.scala 47:24]
  assign _GEN_340 = _T_536 ? _GEN_84 : mem_83; // @[AsyncQueue.scala 47:24]
  assign _GEN_341 = _T_536 ? _GEN_85 : mem_84; // @[AsyncQueue.scala 47:24]
  assign _GEN_342 = _T_536 ? _GEN_86 : mem_85; // @[AsyncQueue.scala 47:24]
  assign _GEN_343 = _T_536 ? _GEN_87 : mem_86; // @[AsyncQueue.scala 47:24]
  assign _GEN_344 = _T_536 ? _GEN_88 : mem_87; // @[AsyncQueue.scala 47:24]
  assign _GEN_345 = _T_536 ? _GEN_89 : mem_88; // @[AsyncQueue.scala 47:24]
  assign _GEN_346 = _T_536 ? _GEN_90 : mem_89; // @[AsyncQueue.scala 47:24]
  assign _GEN_347 = _T_536 ? _GEN_91 : mem_90; // @[AsyncQueue.scala 47:24]
  assign _GEN_348 = _T_536 ? _GEN_92 : mem_91; // @[AsyncQueue.scala 47:24]
  assign _GEN_349 = _T_536 ? _GEN_93 : mem_92; // @[AsyncQueue.scala 47:24]
  assign _GEN_350 = _T_536 ? _GEN_94 : mem_93; // @[AsyncQueue.scala 47:24]
  assign _GEN_351 = _T_536 ? _GEN_95 : mem_94; // @[AsyncQueue.scala 47:24]
  assign _GEN_352 = _T_536 ? _GEN_96 : mem_95; // @[AsyncQueue.scala 47:24]
  assign _GEN_353 = _T_536 ? _GEN_97 : mem_96; // @[AsyncQueue.scala 47:24]
  assign _GEN_354 = _T_536 ? _GEN_98 : mem_97; // @[AsyncQueue.scala 47:24]
  assign _GEN_355 = _T_536 ? _GEN_99 : mem_98; // @[AsyncQueue.scala 47:24]
  assign _GEN_356 = _T_536 ? _GEN_100 : mem_99; // @[AsyncQueue.scala 47:24]
  assign _GEN_357 = _T_536 ? _GEN_101 : mem_100; // @[AsyncQueue.scala 47:24]
  assign _GEN_358 = _T_536 ? _GEN_102 : mem_101; // @[AsyncQueue.scala 47:24]
  assign _GEN_359 = _T_536 ? _GEN_103 : mem_102; // @[AsyncQueue.scala 47:24]
  assign _GEN_360 = _T_536 ? _GEN_104 : mem_103; // @[AsyncQueue.scala 47:24]
  assign _GEN_361 = _T_536 ? _GEN_105 : mem_104; // @[AsyncQueue.scala 47:24]
  assign _GEN_362 = _T_536 ? _GEN_106 : mem_105; // @[AsyncQueue.scala 47:24]
  assign _GEN_363 = _T_536 ? _GEN_107 : mem_106; // @[AsyncQueue.scala 47:24]
  assign _GEN_364 = _T_536 ? _GEN_108 : mem_107; // @[AsyncQueue.scala 47:24]
  assign _GEN_365 = _T_536 ? _GEN_109 : mem_108; // @[AsyncQueue.scala 47:24]
  assign _GEN_366 = _T_536 ? _GEN_110 : mem_109; // @[AsyncQueue.scala 47:24]
  assign _GEN_367 = _T_536 ? _GEN_111 : mem_110; // @[AsyncQueue.scala 47:24]
  assign _GEN_368 = _T_536 ? _GEN_112 : mem_111; // @[AsyncQueue.scala 47:24]
  assign _GEN_369 = _T_536 ? _GEN_113 : mem_112; // @[AsyncQueue.scala 47:24]
  assign _GEN_370 = _T_536 ? _GEN_114 : mem_113; // @[AsyncQueue.scala 47:24]
  assign _GEN_371 = _T_536 ? _GEN_115 : mem_114; // @[AsyncQueue.scala 47:24]
  assign _GEN_372 = _T_536 ? _GEN_116 : mem_115; // @[AsyncQueue.scala 47:24]
  assign _GEN_373 = _T_536 ? _GEN_117 : mem_116; // @[AsyncQueue.scala 47:24]
  assign _GEN_374 = _T_536 ? _GEN_118 : mem_117; // @[AsyncQueue.scala 47:24]
  assign _GEN_375 = _T_536 ? _GEN_119 : mem_118; // @[AsyncQueue.scala 47:24]
  assign _GEN_376 = _T_536 ? _GEN_120 : mem_119; // @[AsyncQueue.scala 47:24]
  assign _GEN_377 = _T_536 ? _GEN_121 : mem_120; // @[AsyncQueue.scala 47:24]
  assign _GEN_378 = _T_536 ? _GEN_122 : mem_121; // @[AsyncQueue.scala 47:24]
  assign _GEN_379 = _T_536 ? _GEN_123 : mem_122; // @[AsyncQueue.scala 47:24]
  assign _GEN_380 = _T_536 ? _GEN_124 : mem_123; // @[AsyncQueue.scala 47:24]
  assign _GEN_381 = _T_536 ? _GEN_125 : mem_124; // @[AsyncQueue.scala 47:24]
  assign _GEN_382 = _T_536 ? _GEN_126 : mem_125; // @[AsyncQueue.scala 47:24]
  assign _GEN_383 = _T_536 ? _GEN_127 : mem_126; // @[AsyncQueue.scala 47:24]
  assign _GEN_384 = _T_536 ? _GEN_128 : mem_127; // @[AsyncQueue.scala 47:24]
  assign _GEN_385 = _T_536 ? _GEN_129 : mem_128; // @[AsyncQueue.scala 47:24]
  assign _GEN_386 = _T_536 ? _GEN_130 : mem_129; // @[AsyncQueue.scala 47:24]
  assign _GEN_387 = _T_536 ? _GEN_131 : mem_130; // @[AsyncQueue.scala 47:24]
  assign _GEN_388 = _T_536 ? _GEN_132 : mem_131; // @[AsyncQueue.scala 47:24]
  assign _GEN_389 = _T_536 ? _GEN_133 : mem_132; // @[AsyncQueue.scala 47:24]
  assign _GEN_390 = _T_536 ? _GEN_134 : mem_133; // @[AsyncQueue.scala 47:24]
  assign _GEN_391 = _T_536 ? _GEN_135 : mem_134; // @[AsyncQueue.scala 47:24]
  assign _GEN_392 = _T_536 ? _GEN_136 : mem_135; // @[AsyncQueue.scala 47:24]
  assign _GEN_393 = _T_536 ? _GEN_137 : mem_136; // @[AsyncQueue.scala 47:24]
  assign _GEN_394 = _T_536 ? _GEN_138 : mem_137; // @[AsyncQueue.scala 47:24]
  assign _GEN_395 = _T_536 ? _GEN_139 : mem_138; // @[AsyncQueue.scala 47:24]
  assign _GEN_396 = _T_536 ? _GEN_140 : mem_139; // @[AsyncQueue.scala 47:24]
  assign _GEN_397 = _T_536 ? _GEN_141 : mem_140; // @[AsyncQueue.scala 47:24]
  assign _GEN_398 = _T_536 ? _GEN_142 : mem_141; // @[AsyncQueue.scala 47:24]
  assign _GEN_399 = _T_536 ? _GEN_143 : mem_142; // @[AsyncQueue.scala 47:24]
  assign _GEN_400 = _T_536 ? _GEN_144 : mem_143; // @[AsyncQueue.scala 47:24]
  assign _GEN_401 = _T_536 ? _GEN_145 : mem_144; // @[AsyncQueue.scala 47:24]
  assign _GEN_402 = _T_536 ? _GEN_146 : mem_145; // @[AsyncQueue.scala 47:24]
  assign _GEN_403 = _T_536 ? _GEN_147 : mem_146; // @[AsyncQueue.scala 47:24]
  assign _GEN_404 = _T_536 ? _GEN_148 : mem_147; // @[AsyncQueue.scala 47:24]
  assign _GEN_405 = _T_536 ? _GEN_149 : mem_148; // @[AsyncQueue.scala 47:24]
  assign _GEN_406 = _T_536 ? _GEN_150 : mem_149; // @[AsyncQueue.scala 47:24]
  assign _GEN_407 = _T_536 ? _GEN_151 : mem_150; // @[AsyncQueue.scala 47:24]
  assign _GEN_408 = _T_536 ? _GEN_152 : mem_151; // @[AsyncQueue.scala 47:24]
  assign _GEN_409 = _T_536 ? _GEN_153 : mem_152; // @[AsyncQueue.scala 47:24]
  assign _GEN_410 = _T_536 ? _GEN_154 : mem_153; // @[AsyncQueue.scala 47:24]
  assign _GEN_411 = _T_536 ? _GEN_155 : mem_154; // @[AsyncQueue.scala 47:24]
  assign _GEN_412 = _T_536 ? _GEN_156 : mem_155; // @[AsyncQueue.scala 47:24]
  assign _GEN_413 = _T_536 ? _GEN_157 : mem_156; // @[AsyncQueue.scala 47:24]
  assign _GEN_414 = _T_536 ? _GEN_158 : mem_157; // @[AsyncQueue.scala 47:24]
  assign _GEN_415 = _T_536 ? _GEN_159 : mem_158; // @[AsyncQueue.scala 47:24]
  assign _GEN_416 = _T_536 ? _GEN_160 : mem_159; // @[AsyncQueue.scala 47:24]
  assign _GEN_417 = _T_536 ? _GEN_161 : mem_160; // @[AsyncQueue.scala 47:24]
  assign _GEN_418 = _T_536 ? _GEN_162 : mem_161; // @[AsyncQueue.scala 47:24]
  assign _GEN_419 = _T_536 ? _GEN_163 : mem_162; // @[AsyncQueue.scala 47:24]
  assign _GEN_420 = _T_536 ? _GEN_164 : mem_163; // @[AsyncQueue.scala 47:24]
  assign _GEN_421 = _T_536 ? _GEN_165 : mem_164; // @[AsyncQueue.scala 47:24]
  assign _GEN_422 = _T_536 ? _GEN_166 : mem_165; // @[AsyncQueue.scala 47:24]
  assign _GEN_423 = _T_536 ? _GEN_167 : mem_166; // @[AsyncQueue.scala 47:24]
  assign _GEN_424 = _T_536 ? _GEN_168 : mem_167; // @[AsyncQueue.scala 47:24]
  assign _GEN_425 = _T_536 ? _GEN_169 : mem_168; // @[AsyncQueue.scala 47:24]
  assign _GEN_426 = _T_536 ? _GEN_170 : mem_169; // @[AsyncQueue.scala 47:24]
  assign _GEN_427 = _T_536 ? _GEN_171 : mem_170; // @[AsyncQueue.scala 47:24]
  assign _GEN_428 = _T_536 ? _GEN_172 : mem_171; // @[AsyncQueue.scala 47:24]
  assign _GEN_429 = _T_536 ? _GEN_173 : mem_172; // @[AsyncQueue.scala 47:24]
  assign _GEN_430 = _T_536 ? _GEN_174 : mem_173; // @[AsyncQueue.scala 47:24]
  assign _GEN_431 = _T_536 ? _GEN_175 : mem_174; // @[AsyncQueue.scala 47:24]
  assign _GEN_432 = _T_536 ? _GEN_176 : mem_175; // @[AsyncQueue.scala 47:24]
  assign _GEN_433 = _T_536 ? _GEN_177 : mem_176; // @[AsyncQueue.scala 47:24]
  assign _GEN_434 = _T_536 ? _GEN_178 : mem_177; // @[AsyncQueue.scala 47:24]
  assign _GEN_435 = _T_536 ? _GEN_179 : mem_178; // @[AsyncQueue.scala 47:24]
  assign _GEN_436 = _T_536 ? _GEN_180 : mem_179; // @[AsyncQueue.scala 47:24]
  assign _GEN_437 = _T_536 ? _GEN_181 : mem_180; // @[AsyncQueue.scala 47:24]
  assign _GEN_438 = _T_536 ? _GEN_182 : mem_181; // @[AsyncQueue.scala 47:24]
  assign _GEN_439 = _T_536 ? _GEN_183 : mem_182; // @[AsyncQueue.scala 47:24]
  assign _GEN_440 = _T_536 ? _GEN_184 : mem_183; // @[AsyncQueue.scala 47:24]
  assign _GEN_441 = _T_536 ? _GEN_185 : mem_184; // @[AsyncQueue.scala 47:24]
  assign _GEN_442 = _T_536 ? _GEN_186 : mem_185; // @[AsyncQueue.scala 47:24]
  assign _GEN_443 = _T_536 ? _GEN_187 : mem_186; // @[AsyncQueue.scala 47:24]
  assign _GEN_444 = _T_536 ? _GEN_188 : mem_187; // @[AsyncQueue.scala 47:24]
  assign _GEN_445 = _T_536 ? _GEN_189 : mem_188; // @[AsyncQueue.scala 47:24]
  assign _GEN_446 = _T_536 ? _GEN_190 : mem_189; // @[AsyncQueue.scala 47:24]
  assign _GEN_447 = _T_536 ? _GEN_191 : mem_190; // @[AsyncQueue.scala 47:24]
  assign _GEN_448 = _T_536 ? _GEN_192 : mem_191; // @[AsyncQueue.scala 47:24]
  assign _GEN_449 = _T_536 ? _GEN_193 : mem_192; // @[AsyncQueue.scala 47:24]
  assign _GEN_450 = _T_536 ? _GEN_194 : mem_193; // @[AsyncQueue.scala 47:24]
  assign _GEN_451 = _T_536 ? _GEN_195 : mem_194; // @[AsyncQueue.scala 47:24]
  assign _GEN_452 = _T_536 ? _GEN_196 : mem_195; // @[AsyncQueue.scala 47:24]
  assign _GEN_453 = _T_536 ? _GEN_197 : mem_196; // @[AsyncQueue.scala 47:24]
  assign _GEN_454 = _T_536 ? _GEN_198 : mem_197; // @[AsyncQueue.scala 47:24]
  assign _GEN_455 = _T_536 ? _GEN_199 : mem_198; // @[AsyncQueue.scala 47:24]
  assign _GEN_456 = _T_536 ? _GEN_200 : mem_199; // @[AsyncQueue.scala 47:24]
  assign _GEN_457 = _T_536 ? _GEN_201 : mem_200; // @[AsyncQueue.scala 47:24]
  assign _GEN_458 = _T_536 ? _GEN_202 : mem_201; // @[AsyncQueue.scala 47:24]
  assign _GEN_459 = _T_536 ? _GEN_203 : mem_202; // @[AsyncQueue.scala 47:24]
  assign _GEN_460 = _T_536 ? _GEN_204 : mem_203; // @[AsyncQueue.scala 47:24]
  assign _GEN_461 = _T_536 ? _GEN_205 : mem_204; // @[AsyncQueue.scala 47:24]
  assign _GEN_462 = _T_536 ? _GEN_206 : mem_205; // @[AsyncQueue.scala 47:24]
  assign _GEN_463 = _T_536 ? _GEN_207 : mem_206; // @[AsyncQueue.scala 47:24]
  assign _GEN_464 = _T_536 ? _GEN_208 : mem_207; // @[AsyncQueue.scala 47:24]
  assign _GEN_465 = _T_536 ? _GEN_209 : mem_208; // @[AsyncQueue.scala 47:24]
  assign _GEN_466 = _T_536 ? _GEN_210 : mem_209; // @[AsyncQueue.scala 47:24]
  assign _GEN_467 = _T_536 ? _GEN_211 : mem_210; // @[AsyncQueue.scala 47:24]
  assign _GEN_468 = _T_536 ? _GEN_212 : mem_211; // @[AsyncQueue.scala 47:24]
  assign _GEN_469 = _T_536 ? _GEN_213 : mem_212; // @[AsyncQueue.scala 47:24]
  assign _GEN_470 = _T_536 ? _GEN_214 : mem_213; // @[AsyncQueue.scala 47:24]
  assign _GEN_471 = _T_536 ? _GEN_215 : mem_214; // @[AsyncQueue.scala 47:24]
  assign _GEN_472 = _T_536 ? _GEN_216 : mem_215; // @[AsyncQueue.scala 47:24]
  assign _GEN_473 = _T_536 ? _GEN_217 : mem_216; // @[AsyncQueue.scala 47:24]
  assign _GEN_474 = _T_536 ? _GEN_218 : mem_217; // @[AsyncQueue.scala 47:24]
  assign _GEN_475 = _T_536 ? _GEN_219 : mem_218; // @[AsyncQueue.scala 47:24]
  assign _GEN_476 = _T_536 ? _GEN_220 : mem_219; // @[AsyncQueue.scala 47:24]
  assign _GEN_477 = _T_536 ? _GEN_221 : mem_220; // @[AsyncQueue.scala 47:24]
  assign _GEN_478 = _T_536 ? _GEN_222 : mem_221; // @[AsyncQueue.scala 47:24]
  assign _GEN_479 = _T_536 ? _GEN_223 : mem_222; // @[AsyncQueue.scala 47:24]
  assign _GEN_480 = _T_536 ? _GEN_224 : mem_223; // @[AsyncQueue.scala 47:24]
  assign _GEN_481 = _T_536 ? _GEN_225 : mem_224; // @[AsyncQueue.scala 47:24]
  assign _GEN_482 = _T_536 ? _GEN_226 : mem_225; // @[AsyncQueue.scala 47:24]
  assign _GEN_483 = _T_536 ? _GEN_227 : mem_226; // @[AsyncQueue.scala 47:24]
  assign _GEN_484 = _T_536 ? _GEN_228 : mem_227; // @[AsyncQueue.scala 47:24]
  assign _GEN_485 = _T_536 ? _GEN_229 : mem_228; // @[AsyncQueue.scala 47:24]
  assign _GEN_486 = _T_536 ? _GEN_230 : mem_229; // @[AsyncQueue.scala 47:24]
  assign _GEN_487 = _T_536 ? _GEN_231 : mem_230; // @[AsyncQueue.scala 47:24]
  assign _GEN_488 = _T_536 ? _GEN_232 : mem_231; // @[AsyncQueue.scala 47:24]
  assign _GEN_489 = _T_536 ? _GEN_233 : mem_232; // @[AsyncQueue.scala 47:24]
  assign _GEN_490 = _T_536 ? _GEN_234 : mem_233; // @[AsyncQueue.scala 47:24]
  assign _GEN_491 = _T_536 ? _GEN_235 : mem_234; // @[AsyncQueue.scala 47:24]
  assign _GEN_492 = _T_536 ? _GEN_236 : mem_235; // @[AsyncQueue.scala 47:24]
  assign _GEN_493 = _T_536 ? _GEN_237 : mem_236; // @[AsyncQueue.scala 47:24]
  assign _GEN_494 = _T_536 ? _GEN_238 : mem_237; // @[AsyncQueue.scala 47:24]
  assign _GEN_495 = _T_536 ? _GEN_239 : mem_238; // @[AsyncQueue.scala 47:24]
  assign _GEN_496 = _T_536 ? _GEN_240 : mem_239; // @[AsyncQueue.scala 47:24]
  assign _GEN_497 = _T_536 ? _GEN_241 : mem_240; // @[AsyncQueue.scala 47:24]
  assign _GEN_498 = _T_536 ? _GEN_242 : mem_241; // @[AsyncQueue.scala 47:24]
  assign _GEN_499 = _T_536 ? _GEN_243 : mem_242; // @[AsyncQueue.scala 47:24]
  assign _GEN_500 = _T_536 ? _GEN_244 : mem_243; // @[AsyncQueue.scala 47:24]
  assign _GEN_501 = _T_536 ? _GEN_245 : mem_244; // @[AsyncQueue.scala 47:24]
  assign _GEN_502 = _T_536 ? _GEN_246 : mem_245; // @[AsyncQueue.scala 47:24]
  assign _GEN_503 = _T_536 ? _GEN_247 : mem_246; // @[AsyncQueue.scala 47:24]
  assign _GEN_504 = _T_536 ? _GEN_248 : mem_247; // @[AsyncQueue.scala 47:24]
  assign _GEN_505 = _T_536 ? _GEN_249 : mem_248; // @[AsyncQueue.scala 47:24]
  assign _GEN_506 = _T_536 ? _GEN_250 : mem_249; // @[AsyncQueue.scala 47:24]
  assign _GEN_507 = _T_536 ? _GEN_251 : mem_250; // @[AsyncQueue.scala 47:24]
  assign _GEN_508 = _T_536 ? _GEN_252 : mem_251; // @[AsyncQueue.scala 47:24]
  assign _GEN_509 = _T_536 ? _GEN_253 : mem_252; // @[AsyncQueue.scala 47:24]
  assign _GEN_510 = _T_536 ? _GEN_254 : mem_253; // @[AsyncQueue.scala 47:24]
  assign _GEN_511 = _T_536 ? _GEN_255 : mem_254; // @[AsyncQueue.scala 47:24]
  assign _GEN_512 = _T_536 ? _GEN_256 : mem_255; // @[AsyncQueue.scala 47:24]
  assign ready_reg_1 = ready_reg_io_q; // @[AsyncQueue.scala 49:59]
  assign _T_558 = ready_reg_1 & sink_ready; // @[AsyncQueue.scala 50:29]
  assign _T_563 = io_sink_reset_n == 1'h0; // @[AsyncQueue.scala 62:36]
  assign _T_564 = reset | _T_563; // @[AsyncQueue.scala 62:33]
  assign io_enq_ready = _T_558;
  assign io_widx = widx_gray_io_q;
  assign io_mem_0 = mem_0;
  assign io_mem_1 = mem_1;
  assign io_mem_2 = mem_2;
  assign io_mem_3 = mem_3;
  assign io_mem_4 = mem_4;
  assign io_mem_5 = mem_5;
  assign io_mem_6 = mem_6;
  assign io_mem_7 = mem_7;
  assign io_mem_8 = mem_8;
  assign io_mem_9 = mem_9;
  assign io_mem_10 = mem_10;
  assign io_mem_11 = mem_11;
  assign io_mem_12 = mem_12;
  assign io_mem_13 = mem_13;
  assign io_mem_14 = mem_14;
  assign io_mem_15 = mem_15;
  assign io_mem_16 = mem_16;
  assign io_mem_17 = mem_17;
  assign io_mem_18 = mem_18;
  assign io_mem_19 = mem_19;
  assign io_mem_20 = mem_20;
  assign io_mem_21 = mem_21;
  assign io_mem_22 = mem_22;
  assign io_mem_23 = mem_23;
  assign io_mem_24 = mem_24;
  assign io_mem_25 = mem_25;
  assign io_mem_26 = mem_26;
  assign io_mem_27 = mem_27;
  assign io_mem_28 = mem_28;
  assign io_mem_29 = mem_29;
  assign io_mem_30 = mem_30;
  assign io_mem_31 = mem_31;
  assign io_mem_32 = mem_32;
  assign io_mem_33 = mem_33;
  assign io_mem_34 = mem_34;
  assign io_mem_35 = mem_35;
  assign io_mem_36 = mem_36;
  assign io_mem_37 = mem_37;
  assign io_mem_38 = mem_38;
  assign io_mem_39 = mem_39;
  assign io_mem_40 = mem_40;
  assign io_mem_41 = mem_41;
  assign io_mem_42 = mem_42;
  assign io_mem_43 = mem_43;
  assign io_mem_44 = mem_44;
  assign io_mem_45 = mem_45;
  assign io_mem_46 = mem_46;
  assign io_mem_47 = mem_47;
  assign io_mem_48 = mem_48;
  assign io_mem_49 = mem_49;
  assign io_mem_50 = mem_50;
  assign io_mem_51 = mem_51;
  assign io_mem_52 = mem_52;
  assign io_mem_53 = mem_53;
  assign io_mem_54 = mem_54;
  assign io_mem_55 = mem_55;
  assign io_mem_56 = mem_56;
  assign io_mem_57 = mem_57;
  assign io_mem_58 = mem_58;
  assign io_mem_59 = mem_59;
  assign io_mem_60 = mem_60;
  assign io_mem_61 = mem_61;
  assign io_mem_62 = mem_62;
  assign io_mem_63 = mem_63;
  assign io_mem_64 = mem_64;
  assign io_mem_65 = mem_65;
  assign io_mem_66 = mem_66;
  assign io_mem_67 = mem_67;
  assign io_mem_68 = mem_68;
  assign io_mem_69 = mem_69;
  assign io_mem_70 = mem_70;
  assign io_mem_71 = mem_71;
  assign io_mem_72 = mem_72;
  assign io_mem_73 = mem_73;
  assign io_mem_74 = mem_74;
  assign io_mem_75 = mem_75;
  assign io_mem_76 = mem_76;
  assign io_mem_77 = mem_77;
  assign io_mem_78 = mem_78;
  assign io_mem_79 = mem_79;
  assign io_mem_80 = mem_80;
  assign io_mem_81 = mem_81;
  assign io_mem_82 = mem_82;
  assign io_mem_83 = mem_83;
  assign io_mem_84 = mem_84;
  assign io_mem_85 = mem_85;
  assign io_mem_86 = mem_86;
  assign io_mem_87 = mem_87;
  assign io_mem_88 = mem_88;
  assign io_mem_89 = mem_89;
  assign io_mem_90 = mem_90;
  assign io_mem_91 = mem_91;
  assign io_mem_92 = mem_92;
  assign io_mem_93 = mem_93;
  assign io_mem_94 = mem_94;
  assign io_mem_95 = mem_95;
  assign io_mem_96 = mem_96;
  assign io_mem_97 = mem_97;
  assign io_mem_98 = mem_98;
  assign io_mem_99 = mem_99;
  assign io_mem_100 = mem_100;
  assign io_mem_101 = mem_101;
  assign io_mem_102 = mem_102;
  assign io_mem_103 = mem_103;
  assign io_mem_104 = mem_104;
  assign io_mem_105 = mem_105;
  assign io_mem_106 = mem_106;
  assign io_mem_107 = mem_107;
  assign io_mem_108 = mem_108;
  assign io_mem_109 = mem_109;
  assign io_mem_110 = mem_110;
  assign io_mem_111 = mem_111;
  assign io_mem_112 = mem_112;
  assign io_mem_113 = mem_113;
  assign io_mem_114 = mem_114;
  assign io_mem_115 = mem_115;
  assign io_mem_116 = mem_116;
  assign io_mem_117 = mem_117;
  assign io_mem_118 = mem_118;
  assign io_mem_119 = mem_119;
  assign io_mem_120 = mem_120;
  assign io_mem_121 = mem_121;
  assign io_mem_122 = mem_122;
  assign io_mem_123 = mem_123;
  assign io_mem_124 = mem_124;
  assign io_mem_125 = mem_125;
  assign io_mem_126 = mem_126;
  assign io_mem_127 = mem_127;
  assign io_mem_128 = mem_128;
  assign io_mem_129 = mem_129;
  assign io_mem_130 = mem_130;
  assign io_mem_131 = mem_131;
  assign io_mem_132 = mem_132;
  assign io_mem_133 = mem_133;
  assign io_mem_134 = mem_134;
  assign io_mem_135 = mem_135;
  assign io_mem_136 = mem_136;
  assign io_mem_137 = mem_137;
  assign io_mem_138 = mem_138;
  assign io_mem_139 = mem_139;
  assign io_mem_140 = mem_140;
  assign io_mem_141 = mem_141;
  assign io_mem_142 = mem_142;
  assign io_mem_143 = mem_143;
  assign io_mem_144 = mem_144;
  assign io_mem_145 = mem_145;
  assign io_mem_146 = mem_146;
  assign io_mem_147 = mem_147;
  assign io_mem_148 = mem_148;
  assign io_mem_149 = mem_149;
  assign io_mem_150 = mem_150;
  assign io_mem_151 = mem_151;
  assign io_mem_152 = mem_152;
  assign io_mem_153 = mem_153;
  assign io_mem_154 = mem_154;
  assign io_mem_155 = mem_155;
  assign io_mem_156 = mem_156;
  assign io_mem_157 = mem_157;
  assign io_mem_158 = mem_158;
  assign io_mem_159 = mem_159;
  assign io_mem_160 = mem_160;
  assign io_mem_161 = mem_161;
  assign io_mem_162 = mem_162;
  assign io_mem_163 = mem_163;
  assign io_mem_164 = mem_164;
  assign io_mem_165 = mem_165;
  assign io_mem_166 = mem_166;
  assign io_mem_167 = mem_167;
  assign io_mem_168 = mem_168;
  assign io_mem_169 = mem_169;
  assign io_mem_170 = mem_170;
  assign io_mem_171 = mem_171;
  assign io_mem_172 = mem_172;
  assign io_mem_173 = mem_173;
  assign io_mem_174 = mem_174;
  assign io_mem_175 = mem_175;
  assign io_mem_176 = mem_176;
  assign io_mem_177 = mem_177;
  assign io_mem_178 = mem_178;
  assign io_mem_179 = mem_179;
  assign io_mem_180 = mem_180;
  assign io_mem_181 = mem_181;
  assign io_mem_182 = mem_182;
  assign io_mem_183 = mem_183;
  assign io_mem_184 = mem_184;
  assign io_mem_185 = mem_185;
  assign io_mem_186 = mem_186;
  assign io_mem_187 = mem_187;
  assign io_mem_188 = mem_188;
  assign io_mem_189 = mem_189;
  assign io_mem_190 = mem_190;
  assign io_mem_191 = mem_191;
  assign io_mem_192 = mem_192;
  assign io_mem_193 = mem_193;
  assign io_mem_194 = mem_194;
  assign io_mem_195 = mem_195;
  assign io_mem_196 = mem_196;
  assign io_mem_197 = mem_197;
  assign io_mem_198 = mem_198;
  assign io_mem_199 = mem_199;
  assign io_mem_200 = mem_200;
  assign io_mem_201 = mem_201;
  assign io_mem_202 = mem_202;
  assign io_mem_203 = mem_203;
  assign io_mem_204 = mem_204;
  assign io_mem_205 = mem_205;
  assign io_mem_206 = mem_206;
  assign io_mem_207 = mem_207;
  assign io_mem_208 = mem_208;
  assign io_mem_209 = mem_209;
  assign io_mem_210 = mem_210;
  assign io_mem_211 = mem_211;
  assign io_mem_212 = mem_212;
  assign io_mem_213 = mem_213;
  assign io_mem_214 = mem_214;
  assign io_mem_215 = mem_215;
  assign io_mem_216 = mem_216;
  assign io_mem_217 = mem_217;
  assign io_mem_218 = mem_218;
  assign io_mem_219 = mem_219;
  assign io_mem_220 = mem_220;
  assign io_mem_221 = mem_221;
  assign io_mem_222 = mem_222;
  assign io_mem_223 = mem_223;
  assign io_mem_224 = mem_224;
  assign io_mem_225 = mem_225;
  assign io_mem_226 = mem_226;
  assign io_mem_227 = mem_227;
  assign io_mem_228 = mem_228;
  assign io_mem_229 = mem_229;
  assign io_mem_230 = mem_230;
  assign io_mem_231 = mem_231;
  assign io_mem_232 = mem_232;
  assign io_mem_233 = mem_233;
  assign io_mem_234 = mem_234;
  assign io_mem_235 = mem_235;
  assign io_mem_236 = mem_236;
  assign io_mem_237 = mem_237;
  assign io_mem_238 = mem_238;
  assign io_mem_239 = mem_239;
  assign io_mem_240 = mem_240;
  assign io_mem_241 = mem_241;
  assign io_mem_242 = mem_242;
  assign io_mem_243 = mem_243;
  assign io_mem_244 = mem_244;
  assign io_mem_245 = mem_245;
  assign io_mem_246 = mem_246;
  assign io_mem_247 = mem_247;
  assign io_mem_248 = mem_248;
  assign io_mem_249 = mem_249;
  assign io_mem_250 = mem_250;
  assign io_mem_251 = mem_251;
  assign io_mem_252 = mem_252;
  assign io_mem_253 = mem_253;
  assign io_mem_254 = mem_254;
  assign io_mem_255 = mem_255;
  assign io_widx_valid = AsyncValidSync_io_out;
  assign widx_bin_clock = clock;
  assign widx_bin_reset = reset;
  assign widx_bin_io_d = _T_545;
  assign widx_bin_io_en = 1'h1;
  assign ridx_gray_clock = clock;
  assign ridx_gray_reset = reset;
  assign ridx_gray_io_d = io_ridx;
  assign ready_reg_clock = clock;
  assign ready_reg_reset = reset;
  assign ready_reg_io_d = ready;
  assign ready_reg_io_en = 1'h1;
  assign widx_gray_clock = clock;
  assign widx_gray_reset = reset;
  assign widx_gray_io_d = widx;
  assign widx_gray_io_en = 1'h1;
  assign AsyncValidSync_clock = clock;
  assign AsyncValidSync_reset = _T_564;
  assign AsyncValidSync_1_clock = clock;
  assign AsyncValidSync_1_reset = _T_564;
  assign AsyncValidSync_1_io_in = io_ridx_valid;
  assign AsyncValidSync_2_clock = clock;
  assign AsyncValidSync_2_reset = reset;
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  mem_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  mem_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  mem_3 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  mem_4 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  mem_5 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  mem_6 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  mem_7 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  mem_8 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  mem_9 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  mem_10 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  mem_11 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  mem_12 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  mem_13 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  mem_14 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  mem_15 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  mem_16 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  mem_17 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  mem_18 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  mem_19 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  mem_20 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  mem_21 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  mem_22 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  mem_23 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  mem_24 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  mem_25 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  mem_26 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  mem_27 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  mem_28 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  mem_29 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  mem_30 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  mem_31 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  mem_32 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  mem_33 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  mem_34 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  mem_35 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  mem_36 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  mem_37 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  mem_38 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  mem_39 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  mem_40 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  mem_41 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  mem_42 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  mem_43 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  mem_44 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  mem_45 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  mem_46 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  mem_47 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  mem_48 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  mem_49 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  mem_50 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  mem_51 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  mem_52 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  mem_53 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  mem_54 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  mem_55 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  mem_56 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  mem_57 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  mem_58 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  mem_59 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  mem_60 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  mem_61 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  mem_62 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  mem_63 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  mem_64 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  mem_65 = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  mem_66 = _RAND_66[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  mem_67 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  mem_68 = _RAND_68[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  mem_69 = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  mem_70 = _RAND_70[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  mem_71 = _RAND_71[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  mem_72 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  mem_73 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  mem_74 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  mem_75 = _RAND_75[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  mem_76 = _RAND_76[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  mem_77 = _RAND_77[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  mem_78 = _RAND_78[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  mem_79 = _RAND_79[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  mem_80 = _RAND_80[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  mem_81 = _RAND_81[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  mem_82 = _RAND_82[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  mem_83 = _RAND_83[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  mem_84 = _RAND_84[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  mem_85 = _RAND_85[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  mem_86 = _RAND_86[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  mem_87 = _RAND_87[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  mem_88 = _RAND_88[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  mem_89 = _RAND_89[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  mem_90 = _RAND_90[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  mem_91 = _RAND_91[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  mem_92 = _RAND_92[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  mem_93 = _RAND_93[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  mem_94 = _RAND_94[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  mem_95 = _RAND_95[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  mem_96 = _RAND_96[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  mem_97 = _RAND_97[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  mem_98 = _RAND_98[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  mem_99 = _RAND_99[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  mem_100 = _RAND_100[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  mem_101 = _RAND_101[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  mem_102 = _RAND_102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  mem_103 = _RAND_103[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  mem_104 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  mem_105 = _RAND_105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  mem_106 = _RAND_106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  mem_107 = _RAND_107[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  mem_108 = _RAND_108[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  mem_109 = _RAND_109[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  mem_110 = _RAND_110[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  mem_111 = _RAND_111[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  mem_112 = _RAND_112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  mem_113 = _RAND_113[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  mem_114 = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  mem_115 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  mem_116 = _RAND_116[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  mem_117 = _RAND_117[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  mem_118 = _RAND_118[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  mem_119 = _RAND_119[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  mem_120 = _RAND_120[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  mem_121 = _RAND_121[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  mem_122 = _RAND_122[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  mem_123 = _RAND_123[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  mem_124 = _RAND_124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  mem_125 = _RAND_125[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  mem_126 = _RAND_126[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  mem_127 = _RAND_127[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  mem_128 = _RAND_128[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  mem_129 = _RAND_129[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  mem_130 = _RAND_130[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  mem_131 = _RAND_131[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  mem_132 = _RAND_132[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  mem_133 = _RAND_133[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  mem_134 = _RAND_134[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  mem_135 = _RAND_135[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  mem_136 = _RAND_136[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  mem_137 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  mem_138 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  mem_139 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  mem_140 = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  mem_141 = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  mem_142 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  mem_143 = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  mem_144 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  mem_145 = _RAND_145[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  mem_146 = _RAND_146[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  mem_147 = _RAND_147[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  mem_148 = _RAND_148[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  mem_149 = _RAND_149[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  mem_150 = _RAND_150[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  mem_151 = _RAND_151[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  mem_152 = _RAND_152[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  mem_153 = _RAND_153[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  mem_154 = _RAND_154[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  mem_155 = _RAND_155[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  mem_156 = _RAND_156[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  mem_157 = _RAND_157[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  mem_158 = _RAND_158[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  mem_159 = _RAND_159[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  mem_160 = _RAND_160[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  mem_161 = _RAND_161[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  mem_162 = _RAND_162[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  mem_163 = _RAND_163[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  mem_164 = _RAND_164[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  mem_165 = _RAND_165[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  mem_166 = _RAND_166[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  mem_167 = _RAND_167[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  mem_168 = _RAND_168[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  mem_169 = _RAND_169[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  mem_170 = _RAND_170[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  mem_171 = _RAND_171[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  mem_172 = _RAND_172[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  mem_173 = _RAND_173[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  mem_174 = _RAND_174[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  mem_175 = _RAND_175[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  mem_176 = _RAND_176[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  mem_177 = _RAND_177[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  mem_178 = _RAND_178[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  mem_179 = _RAND_179[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  mem_180 = _RAND_180[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  mem_181 = _RAND_181[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  mem_182 = _RAND_182[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  mem_183 = _RAND_183[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  mem_184 = _RAND_184[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  mem_185 = _RAND_185[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  mem_186 = _RAND_186[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  mem_187 = _RAND_187[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  mem_188 = _RAND_188[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  mem_189 = _RAND_189[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  mem_190 = _RAND_190[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  mem_191 = _RAND_191[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  mem_192 = _RAND_192[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  mem_193 = _RAND_193[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{$random}};
  mem_194 = _RAND_194[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{$random}};
  mem_195 = _RAND_195[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{$random}};
  mem_196 = _RAND_196[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{$random}};
  mem_197 = _RAND_197[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{$random}};
  mem_198 = _RAND_198[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{$random}};
  mem_199 = _RAND_199[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{$random}};
  mem_200 = _RAND_200[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{$random}};
  mem_201 = _RAND_201[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{$random}};
  mem_202 = _RAND_202[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{$random}};
  mem_203 = _RAND_203[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{$random}};
  mem_204 = _RAND_204[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{$random}};
  mem_205 = _RAND_205[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{$random}};
  mem_206 = _RAND_206[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{$random}};
  mem_207 = _RAND_207[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{$random}};
  mem_208 = _RAND_208[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{$random}};
  mem_209 = _RAND_209[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{$random}};
  mem_210 = _RAND_210[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{$random}};
  mem_211 = _RAND_211[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{$random}};
  mem_212 = _RAND_212[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{$random}};
  mem_213 = _RAND_213[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{$random}};
  mem_214 = _RAND_214[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{$random}};
  mem_215 = _RAND_215[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{$random}};
  mem_216 = _RAND_216[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{$random}};
  mem_217 = _RAND_217[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{$random}};
  mem_218 = _RAND_218[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{$random}};
  mem_219 = _RAND_219[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{$random}};
  mem_220 = _RAND_220[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{$random}};
  mem_221 = _RAND_221[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{$random}};
  mem_222 = _RAND_222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{$random}};
  mem_223 = _RAND_223[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{$random}};
  mem_224 = _RAND_224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{$random}};
  mem_225 = _RAND_225[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{$random}};
  mem_226 = _RAND_226[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{$random}};
  mem_227 = _RAND_227[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{$random}};
  mem_228 = _RAND_228[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{$random}};
  mem_229 = _RAND_229[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{$random}};
  mem_230 = _RAND_230[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{$random}};
  mem_231 = _RAND_231[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{$random}};
  mem_232 = _RAND_232[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{$random}};
  mem_233 = _RAND_233[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{$random}};
  mem_234 = _RAND_234[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{$random}};
  mem_235 = _RAND_235[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{$random}};
  mem_236 = _RAND_236[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{$random}};
  mem_237 = _RAND_237[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{$random}};
  mem_238 = _RAND_238[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{$random}};
  mem_239 = _RAND_239[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{$random}};
  mem_240 = _RAND_240[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{$random}};
  mem_241 = _RAND_241[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{$random}};
  mem_242 = _RAND_242[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{$random}};
  mem_243 = _RAND_243[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{$random}};
  mem_244 = _RAND_244[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{$random}};
  mem_245 = _RAND_245[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{$random}};
  mem_246 = _RAND_246[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{$random}};
  mem_247 = _RAND_247[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{$random}};
  mem_248 = _RAND_248[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{$random}};
  mem_249 = _RAND_249[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{$random}};
  mem_250 = _RAND_250[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{$random}};
  mem_251 = _RAND_251[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{$random}};
  mem_252 = _RAND_252[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{$random}};
  mem_253 = _RAND_253[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{$random}};
  mem_254 = _RAND_254[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{$random}};
  mem_255 = _RAND_255[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_536) begin
      if (8'h0 == index) begin
        mem_0 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1 == index) begin
        mem_1 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2 == index) begin
        mem_2 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3 == index) begin
        mem_3 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4 == index) begin
        mem_4 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5 == index) begin
        mem_5 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6 == index) begin
        mem_6 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7 == index) begin
        mem_7 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8 == index) begin
        mem_8 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9 == index) begin
        mem_9 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha == index) begin
        mem_10 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb == index) begin
        mem_11 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc == index) begin
        mem_12 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd == index) begin
        mem_13 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he == index) begin
        mem_14 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf == index) begin
        mem_15 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h10 == index) begin
        mem_16 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h11 == index) begin
        mem_17 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h12 == index) begin
        mem_18 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h13 == index) begin
        mem_19 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h14 == index) begin
        mem_20 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h15 == index) begin
        mem_21 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h16 == index) begin
        mem_22 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h17 == index) begin
        mem_23 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h18 == index) begin
        mem_24 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h19 == index) begin
        mem_25 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1a == index) begin
        mem_26 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1b == index) begin
        mem_27 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1c == index) begin
        mem_28 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1d == index) begin
        mem_29 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1e == index) begin
        mem_30 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h1f == index) begin
        mem_31 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h20 == index) begin
        mem_32 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h21 == index) begin
        mem_33 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h22 == index) begin
        mem_34 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h23 == index) begin
        mem_35 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h24 == index) begin
        mem_36 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h25 == index) begin
        mem_37 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h26 == index) begin
        mem_38 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h27 == index) begin
        mem_39 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h28 == index) begin
        mem_40 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h29 == index) begin
        mem_41 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2a == index) begin
        mem_42 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2b == index) begin
        mem_43 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2c == index) begin
        mem_44 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2d == index) begin
        mem_45 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2e == index) begin
        mem_46 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h2f == index) begin
        mem_47 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h30 == index) begin
        mem_48 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h31 == index) begin
        mem_49 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h32 == index) begin
        mem_50 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h33 == index) begin
        mem_51 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h34 == index) begin
        mem_52 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h35 == index) begin
        mem_53 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h36 == index) begin
        mem_54 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h37 == index) begin
        mem_55 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h38 == index) begin
        mem_56 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h39 == index) begin
        mem_57 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3a == index) begin
        mem_58 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3b == index) begin
        mem_59 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3c == index) begin
        mem_60 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3d == index) begin
        mem_61 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3e == index) begin
        mem_62 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h3f == index) begin
        mem_63 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h40 == index) begin
        mem_64 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h41 == index) begin
        mem_65 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h42 == index) begin
        mem_66 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h43 == index) begin
        mem_67 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h44 == index) begin
        mem_68 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h45 == index) begin
        mem_69 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h46 == index) begin
        mem_70 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h47 == index) begin
        mem_71 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h48 == index) begin
        mem_72 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h49 == index) begin
        mem_73 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4a == index) begin
        mem_74 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4b == index) begin
        mem_75 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4c == index) begin
        mem_76 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4d == index) begin
        mem_77 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4e == index) begin
        mem_78 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h4f == index) begin
        mem_79 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h50 == index) begin
        mem_80 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h51 == index) begin
        mem_81 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h52 == index) begin
        mem_82 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h53 == index) begin
        mem_83 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h54 == index) begin
        mem_84 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h55 == index) begin
        mem_85 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h56 == index) begin
        mem_86 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h57 == index) begin
        mem_87 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h58 == index) begin
        mem_88 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h59 == index) begin
        mem_89 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5a == index) begin
        mem_90 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5b == index) begin
        mem_91 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5c == index) begin
        mem_92 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5d == index) begin
        mem_93 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5e == index) begin
        mem_94 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h5f == index) begin
        mem_95 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h60 == index) begin
        mem_96 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h61 == index) begin
        mem_97 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h62 == index) begin
        mem_98 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h63 == index) begin
        mem_99 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h64 == index) begin
        mem_100 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h65 == index) begin
        mem_101 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h66 == index) begin
        mem_102 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h67 == index) begin
        mem_103 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h68 == index) begin
        mem_104 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h69 == index) begin
        mem_105 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6a == index) begin
        mem_106 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6b == index) begin
        mem_107 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6c == index) begin
        mem_108 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6d == index) begin
        mem_109 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6e == index) begin
        mem_110 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h6f == index) begin
        mem_111 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h70 == index) begin
        mem_112 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h71 == index) begin
        mem_113 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h72 == index) begin
        mem_114 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h73 == index) begin
        mem_115 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h74 == index) begin
        mem_116 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h75 == index) begin
        mem_117 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h76 == index) begin
        mem_118 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h77 == index) begin
        mem_119 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h78 == index) begin
        mem_120 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h79 == index) begin
        mem_121 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7a == index) begin
        mem_122 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7b == index) begin
        mem_123 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7c == index) begin
        mem_124 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7d == index) begin
        mem_125 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7e == index) begin
        mem_126 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h7f == index) begin
        mem_127 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h80 == index) begin
        mem_128 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h81 == index) begin
        mem_129 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h82 == index) begin
        mem_130 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h83 == index) begin
        mem_131 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h84 == index) begin
        mem_132 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h85 == index) begin
        mem_133 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h86 == index) begin
        mem_134 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h87 == index) begin
        mem_135 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h88 == index) begin
        mem_136 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h89 == index) begin
        mem_137 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8a == index) begin
        mem_138 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8b == index) begin
        mem_139 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8c == index) begin
        mem_140 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8d == index) begin
        mem_141 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8e == index) begin
        mem_142 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h8f == index) begin
        mem_143 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h90 == index) begin
        mem_144 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h91 == index) begin
        mem_145 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h92 == index) begin
        mem_146 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h93 == index) begin
        mem_147 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h94 == index) begin
        mem_148 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h95 == index) begin
        mem_149 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h96 == index) begin
        mem_150 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h97 == index) begin
        mem_151 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h98 == index) begin
        mem_152 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h99 == index) begin
        mem_153 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9a == index) begin
        mem_154 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9b == index) begin
        mem_155 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9c == index) begin
        mem_156 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9d == index) begin
        mem_157 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9e == index) begin
        mem_158 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'h9f == index) begin
        mem_159 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha0 == index) begin
        mem_160 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha1 == index) begin
        mem_161 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha2 == index) begin
        mem_162 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha3 == index) begin
        mem_163 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha4 == index) begin
        mem_164 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha5 == index) begin
        mem_165 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha6 == index) begin
        mem_166 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha7 == index) begin
        mem_167 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha8 == index) begin
        mem_168 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'ha9 == index) begin
        mem_169 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'haa == index) begin
        mem_170 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hab == index) begin
        mem_171 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hac == index) begin
        mem_172 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'had == index) begin
        mem_173 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hae == index) begin
        mem_174 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'haf == index) begin
        mem_175 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb0 == index) begin
        mem_176 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb1 == index) begin
        mem_177 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb2 == index) begin
        mem_178 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb3 == index) begin
        mem_179 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb4 == index) begin
        mem_180 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb5 == index) begin
        mem_181 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb6 == index) begin
        mem_182 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb7 == index) begin
        mem_183 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb8 == index) begin
        mem_184 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hb9 == index) begin
        mem_185 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hba == index) begin
        mem_186 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hbb == index) begin
        mem_187 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hbc == index) begin
        mem_188 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hbd == index) begin
        mem_189 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hbe == index) begin
        mem_190 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hbf == index) begin
        mem_191 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc0 == index) begin
        mem_192 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc1 == index) begin
        mem_193 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc2 == index) begin
        mem_194 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc3 == index) begin
        mem_195 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc4 == index) begin
        mem_196 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc5 == index) begin
        mem_197 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc6 == index) begin
        mem_198 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc7 == index) begin
        mem_199 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc8 == index) begin
        mem_200 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hc9 == index) begin
        mem_201 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hca == index) begin
        mem_202 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hcb == index) begin
        mem_203 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hcc == index) begin
        mem_204 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hcd == index) begin
        mem_205 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hce == index) begin
        mem_206 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hcf == index) begin
        mem_207 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd0 == index) begin
        mem_208 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd1 == index) begin
        mem_209 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd2 == index) begin
        mem_210 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd3 == index) begin
        mem_211 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd4 == index) begin
        mem_212 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd5 == index) begin
        mem_213 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd6 == index) begin
        mem_214 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd7 == index) begin
        mem_215 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd8 == index) begin
        mem_216 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hd9 == index) begin
        mem_217 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hda == index) begin
        mem_218 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hdb == index) begin
        mem_219 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hdc == index) begin
        mem_220 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hdd == index) begin
        mem_221 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hde == index) begin
        mem_222 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hdf == index) begin
        mem_223 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he0 == index) begin
        mem_224 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he1 == index) begin
        mem_225 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he2 == index) begin
        mem_226 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he3 == index) begin
        mem_227 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he4 == index) begin
        mem_228 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he5 == index) begin
        mem_229 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he6 == index) begin
        mem_230 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he7 == index) begin
        mem_231 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he8 == index) begin
        mem_232 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'he9 == index) begin
        mem_233 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hea == index) begin
        mem_234 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'heb == index) begin
        mem_235 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hec == index) begin
        mem_236 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hed == index) begin
        mem_237 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hee == index) begin
        mem_238 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hef == index) begin
        mem_239 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf0 == index) begin
        mem_240 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf1 == index) begin
        mem_241 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf2 == index) begin
        mem_242 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf3 == index) begin
        mem_243 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf4 == index) begin
        mem_244 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf5 == index) begin
        mem_245 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf6 == index) begin
        mem_246 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf7 == index) begin
        mem_247 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf8 == index) begin
        mem_248 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hf9 == index) begin
        mem_249 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hfa == index) begin
        mem_250 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hfb == index) begin
        mem_251 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hfc == index) begin
        mem_252 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hfd == index) begin
        mem_253 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hfe == index) begin
        mem_254 <= io_enq_bits;
      end
    end
    if (_T_536) begin
      if (8'hff == index) begin
        mem_255 <= io_enq_bits;
      end
    end
  end
endmodule
module SynchronizerShiftReg_w8_d1(
  input        clock,
  input  [7:0] io_d,
  output [7:0] io_q
);
  reg [7:0] sync_0; // @[ShiftReg.scala 114:16]
  reg [31:0] _RAND_0;
  assign io_q = sync_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  sync_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    sync_0 <= io_d;
  end
endmodule
module AsyncQueueSink_1(
  input        clock,
  input        reset,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output [8:0] io_ridx,
  input  [8:0] io_widx,
  input  [7:0] io_mem_0,
  input  [7:0] io_mem_1,
  input  [7:0] io_mem_2,
  input  [7:0] io_mem_3,
  input  [7:0] io_mem_4,
  input  [7:0] io_mem_5,
  input  [7:0] io_mem_6,
  input  [7:0] io_mem_7,
  input  [7:0] io_mem_8,
  input  [7:0] io_mem_9,
  input  [7:0] io_mem_10,
  input  [7:0] io_mem_11,
  input  [7:0] io_mem_12,
  input  [7:0] io_mem_13,
  input  [7:0] io_mem_14,
  input  [7:0] io_mem_15,
  input  [7:0] io_mem_16,
  input  [7:0] io_mem_17,
  input  [7:0] io_mem_18,
  input  [7:0] io_mem_19,
  input  [7:0] io_mem_20,
  input  [7:0] io_mem_21,
  input  [7:0] io_mem_22,
  input  [7:0] io_mem_23,
  input  [7:0] io_mem_24,
  input  [7:0] io_mem_25,
  input  [7:0] io_mem_26,
  input  [7:0] io_mem_27,
  input  [7:0] io_mem_28,
  input  [7:0] io_mem_29,
  input  [7:0] io_mem_30,
  input  [7:0] io_mem_31,
  input  [7:0] io_mem_32,
  input  [7:0] io_mem_33,
  input  [7:0] io_mem_34,
  input  [7:0] io_mem_35,
  input  [7:0] io_mem_36,
  input  [7:0] io_mem_37,
  input  [7:0] io_mem_38,
  input  [7:0] io_mem_39,
  input  [7:0] io_mem_40,
  input  [7:0] io_mem_41,
  input  [7:0] io_mem_42,
  input  [7:0] io_mem_43,
  input  [7:0] io_mem_44,
  input  [7:0] io_mem_45,
  input  [7:0] io_mem_46,
  input  [7:0] io_mem_47,
  input  [7:0] io_mem_48,
  input  [7:0] io_mem_49,
  input  [7:0] io_mem_50,
  input  [7:0] io_mem_51,
  input  [7:0] io_mem_52,
  input  [7:0] io_mem_53,
  input  [7:0] io_mem_54,
  input  [7:0] io_mem_55,
  input  [7:0] io_mem_56,
  input  [7:0] io_mem_57,
  input  [7:0] io_mem_58,
  input  [7:0] io_mem_59,
  input  [7:0] io_mem_60,
  input  [7:0] io_mem_61,
  input  [7:0] io_mem_62,
  input  [7:0] io_mem_63,
  input  [7:0] io_mem_64,
  input  [7:0] io_mem_65,
  input  [7:0] io_mem_66,
  input  [7:0] io_mem_67,
  input  [7:0] io_mem_68,
  input  [7:0] io_mem_69,
  input  [7:0] io_mem_70,
  input  [7:0] io_mem_71,
  input  [7:0] io_mem_72,
  input  [7:0] io_mem_73,
  input  [7:0] io_mem_74,
  input  [7:0] io_mem_75,
  input  [7:0] io_mem_76,
  input  [7:0] io_mem_77,
  input  [7:0] io_mem_78,
  input  [7:0] io_mem_79,
  input  [7:0] io_mem_80,
  input  [7:0] io_mem_81,
  input  [7:0] io_mem_82,
  input  [7:0] io_mem_83,
  input  [7:0] io_mem_84,
  input  [7:0] io_mem_85,
  input  [7:0] io_mem_86,
  input  [7:0] io_mem_87,
  input  [7:0] io_mem_88,
  input  [7:0] io_mem_89,
  input  [7:0] io_mem_90,
  input  [7:0] io_mem_91,
  input  [7:0] io_mem_92,
  input  [7:0] io_mem_93,
  input  [7:0] io_mem_94,
  input  [7:0] io_mem_95,
  input  [7:0] io_mem_96,
  input  [7:0] io_mem_97,
  input  [7:0] io_mem_98,
  input  [7:0] io_mem_99,
  input  [7:0] io_mem_100,
  input  [7:0] io_mem_101,
  input  [7:0] io_mem_102,
  input  [7:0] io_mem_103,
  input  [7:0] io_mem_104,
  input  [7:0] io_mem_105,
  input  [7:0] io_mem_106,
  input  [7:0] io_mem_107,
  input  [7:0] io_mem_108,
  input  [7:0] io_mem_109,
  input  [7:0] io_mem_110,
  input  [7:0] io_mem_111,
  input  [7:0] io_mem_112,
  input  [7:0] io_mem_113,
  input  [7:0] io_mem_114,
  input  [7:0] io_mem_115,
  input  [7:0] io_mem_116,
  input  [7:0] io_mem_117,
  input  [7:0] io_mem_118,
  input  [7:0] io_mem_119,
  input  [7:0] io_mem_120,
  input  [7:0] io_mem_121,
  input  [7:0] io_mem_122,
  input  [7:0] io_mem_123,
  input  [7:0] io_mem_124,
  input  [7:0] io_mem_125,
  input  [7:0] io_mem_126,
  input  [7:0] io_mem_127,
  input  [7:0] io_mem_128,
  input  [7:0] io_mem_129,
  input  [7:0] io_mem_130,
  input  [7:0] io_mem_131,
  input  [7:0] io_mem_132,
  input  [7:0] io_mem_133,
  input  [7:0] io_mem_134,
  input  [7:0] io_mem_135,
  input  [7:0] io_mem_136,
  input  [7:0] io_mem_137,
  input  [7:0] io_mem_138,
  input  [7:0] io_mem_139,
  input  [7:0] io_mem_140,
  input  [7:0] io_mem_141,
  input  [7:0] io_mem_142,
  input  [7:0] io_mem_143,
  input  [7:0] io_mem_144,
  input  [7:0] io_mem_145,
  input  [7:0] io_mem_146,
  input  [7:0] io_mem_147,
  input  [7:0] io_mem_148,
  input  [7:0] io_mem_149,
  input  [7:0] io_mem_150,
  input  [7:0] io_mem_151,
  input  [7:0] io_mem_152,
  input  [7:0] io_mem_153,
  input  [7:0] io_mem_154,
  input  [7:0] io_mem_155,
  input  [7:0] io_mem_156,
  input  [7:0] io_mem_157,
  input  [7:0] io_mem_158,
  input  [7:0] io_mem_159,
  input  [7:0] io_mem_160,
  input  [7:0] io_mem_161,
  input  [7:0] io_mem_162,
  input  [7:0] io_mem_163,
  input  [7:0] io_mem_164,
  input  [7:0] io_mem_165,
  input  [7:0] io_mem_166,
  input  [7:0] io_mem_167,
  input  [7:0] io_mem_168,
  input  [7:0] io_mem_169,
  input  [7:0] io_mem_170,
  input  [7:0] io_mem_171,
  input  [7:0] io_mem_172,
  input  [7:0] io_mem_173,
  input  [7:0] io_mem_174,
  input  [7:0] io_mem_175,
  input  [7:0] io_mem_176,
  input  [7:0] io_mem_177,
  input  [7:0] io_mem_178,
  input  [7:0] io_mem_179,
  input  [7:0] io_mem_180,
  input  [7:0] io_mem_181,
  input  [7:0] io_mem_182,
  input  [7:0] io_mem_183,
  input  [7:0] io_mem_184,
  input  [7:0] io_mem_185,
  input  [7:0] io_mem_186,
  input  [7:0] io_mem_187,
  input  [7:0] io_mem_188,
  input  [7:0] io_mem_189,
  input  [7:0] io_mem_190,
  input  [7:0] io_mem_191,
  input  [7:0] io_mem_192,
  input  [7:0] io_mem_193,
  input  [7:0] io_mem_194,
  input  [7:0] io_mem_195,
  input  [7:0] io_mem_196,
  input  [7:0] io_mem_197,
  input  [7:0] io_mem_198,
  input  [7:0] io_mem_199,
  input  [7:0] io_mem_200,
  input  [7:0] io_mem_201,
  input  [7:0] io_mem_202,
  input  [7:0] io_mem_203,
  input  [7:0] io_mem_204,
  input  [7:0] io_mem_205,
  input  [7:0] io_mem_206,
  input  [7:0] io_mem_207,
  input  [7:0] io_mem_208,
  input  [7:0] io_mem_209,
  input  [7:0] io_mem_210,
  input  [7:0] io_mem_211,
  input  [7:0] io_mem_212,
  input  [7:0] io_mem_213,
  input  [7:0] io_mem_214,
  input  [7:0] io_mem_215,
  input  [7:0] io_mem_216,
  input  [7:0] io_mem_217,
  input  [7:0] io_mem_218,
  input  [7:0] io_mem_219,
  input  [7:0] io_mem_220,
  input  [7:0] io_mem_221,
  input  [7:0] io_mem_222,
  input  [7:0] io_mem_223,
  input  [7:0] io_mem_224,
  input  [7:0] io_mem_225,
  input  [7:0] io_mem_226,
  input  [7:0] io_mem_227,
  input  [7:0] io_mem_228,
  input  [7:0] io_mem_229,
  input  [7:0] io_mem_230,
  input  [7:0] io_mem_231,
  input  [7:0] io_mem_232,
  input  [7:0] io_mem_233,
  input  [7:0] io_mem_234,
  input  [7:0] io_mem_235,
  input  [7:0] io_mem_236,
  input  [7:0] io_mem_237,
  input  [7:0] io_mem_238,
  input  [7:0] io_mem_239,
  input  [7:0] io_mem_240,
  input  [7:0] io_mem_241,
  input  [7:0] io_mem_242,
  input  [7:0] io_mem_243,
  input  [7:0] io_mem_244,
  input  [7:0] io_mem_245,
  input  [7:0] io_mem_246,
  input  [7:0] io_mem_247,
  input  [7:0] io_mem_248,
  input  [7:0] io_mem_249,
  input  [7:0] io_mem_250,
  input  [7:0] io_mem_251,
  input  [7:0] io_mem_252,
  input  [7:0] io_mem_253,
  input  [7:0] io_mem_254,
  input  [7:0] io_mem_255,
  input        io_source_reset_n,
  output       io_ridx_valid,
  input        io_widx_valid
);
  wire  ridx_bin_clock; // @[AsyncResetReg.scala 110:21]
  wire  ridx_bin_reset; // @[AsyncResetReg.scala 110:21]
  wire [8:0] ridx_bin_io_d; // @[AsyncResetReg.scala 110:21]
  wire [8:0] ridx_bin_io_q; // @[AsyncResetReg.scala 110:21]
  wire  ridx_bin_io_en; // @[AsyncResetReg.scala 110:21]
  wire  widx_gray_clock; // @[ShiftReg.scala 47:23]
  wire  widx_gray_reset; // @[ShiftReg.scala 47:23]
  wire [8:0] widx_gray_io_d; // @[ShiftReg.scala 47:23]
  wire [8:0] widx_gray_io_q; // @[ShiftReg.scala 47:23]
  wire  deq_bits_reg_clock; // @[ShiftReg.scala 47:23]
  wire [7:0] deq_bits_reg_io_d; // @[ShiftReg.scala 47:23]
  wire [7:0] deq_bits_reg_io_q; // @[ShiftReg.scala 47:23]
  wire  valid_reg_clock; // @[AsyncResetReg.scala 110:21]
  wire  valid_reg_reset; // @[AsyncResetReg.scala 110:21]
  wire  valid_reg_io_d; // @[AsyncResetReg.scala 110:21]
  wire  valid_reg_io_q; // @[AsyncResetReg.scala 110:21]
  wire  valid_reg_io_en; // @[AsyncResetReg.scala 110:21]
  wire  ridx_gray_clock; // @[AsyncResetReg.scala 110:21]
  wire  ridx_gray_reset; // @[AsyncResetReg.scala 110:21]
  wire [8:0] ridx_gray_io_d; // @[AsyncResetReg.scala 110:21]
  wire [8:0] ridx_gray_io_q; // @[AsyncResetReg.scala 110:21]
  wire  ridx_gray_io_en; // @[AsyncResetReg.scala 110:21]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 124:31]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 124:31]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 124:31]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 125:31]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 125:31]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 125:31]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 125:31]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 126:31]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 126:31]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 126:31]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 126:31]
  wire  AsyncResetRegVec_w1_i0_clock; // @[AsyncResetReg.scala 110:21]
  wire  AsyncResetRegVec_w1_i0_reset; // @[AsyncResetReg.scala 110:21]
  wire  AsyncResetRegVec_w1_i0_io_d; // @[AsyncResetReg.scala 110:21]
  wire  AsyncResetRegVec_w1_i0_io_q; // @[AsyncResetReg.scala 110:21]
  wire  AsyncResetRegVec_w1_i0_io_en; // @[AsyncResetReg.scala 110:21]
  wire  _T_272; // @[Decoupled.scala 30:37]
  wire  source_ready;
  wire  _T_274; // @[AsyncQueue.scala 99:49]
  wire [8:0] _GEN_256; // @[AsyncQueue.scala 11:47]
  wire [9:0] _T_279; // @[AsyncQueue.scala 11:47]
  wire [8:0] _T_280; // @[AsyncQueue.scala 11:47]
  wire [8:0] _T_281; // @[AsyncQueue.scala 11:23]
  wire [8:0] _T_283; // @[AsyncQueue.scala 12:32]
  wire [8:0] ridx; // @[AsyncQueue.scala 12:17]
  wire [8:0] widx; // @[ShiftReg.scala 50:24]
  wire  _T_285; // @[AsyncQueue.scala 101:36]
  wire  valid; // @[AsyncQueue.scala 101:28]
  wire [7:0] _T_286; // @[AsyncQueue.scala 107:48]
  wire  _T_287; // @[AsyncQueue.scala 107:67]
  wire [7:0] _GEN_257; // @[AsyncQueue.scala 107:80]
  wire [7:0] _T_288; // @[AsyncQueue.scala 107:80]
  wire [7:0] index; // @[AsyncQueue.scala 107:60]
  wire [7:0] _GEN_1; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_2; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_3; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_4; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_5; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_6; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_7; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_8; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_9; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_10; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_11; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_12; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_13; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_14; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_15; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_16; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_17; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_18; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_19; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_20; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_21; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_22; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_23; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_24; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_25; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_26; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_27; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_28; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_29; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_30; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_31; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_32; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_33; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_34; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_35; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_36; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_37; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_38; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_39; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_40; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_41; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_42; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_43; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_44; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_45; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_46; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_47; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_48; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_49; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_50; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_51; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_52; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_53; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_54; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_55; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_56; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_57; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_58; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_59; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_60; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_61; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_62; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_63; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_64; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_65; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_66; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_67; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_68; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_69; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_70; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_71; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_72; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_73; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_74; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_75; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_76; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_77; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_78; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_79; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_80; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_81; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_82; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_83; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_84; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_85; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_86; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_87; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_88; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_89; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_90; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_91; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_92; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_93; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_94; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_95; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_96; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_97; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_98; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_99; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_100; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_101; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_102; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_103; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_104; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_105; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_106; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_107; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_108; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_109; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_110; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_111; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_112; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_113; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_114; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_115; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_116; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_117; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_118; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_119; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_120; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_121; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_122; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_123; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_124; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_125; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_126; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_127; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_128; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_129; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_130; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_131; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_132; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_133; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_134; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_135; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_136; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_137; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_138; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_139; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_140; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_141; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_142; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_143; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_144; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_145; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_146; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_147; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_148; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_149; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_150; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_151; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_152; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_153; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_154; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_155; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_156; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_157; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_158; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_159; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_160; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_161; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_162; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_163; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_164; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_165; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_166; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_167; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_168; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_169; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_170; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_171; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_172; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_173; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_174; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_175; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_176; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_177; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_178; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_179; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_180; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_181; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_182; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_183; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_184; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_185; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_186; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_187; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_188; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_189; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_190; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_191; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_192; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_193; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_194; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_195; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_196; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_197; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_198; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_199; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_200; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_201; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_202; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_203; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_204; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_205; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_206; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_207; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_208; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_209; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_210; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_211; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_212; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_213; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_214; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_215; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_216; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_217; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_218; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_219; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_220; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_221; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_222; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_223; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_224; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_225; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_226; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_227; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_228; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_229; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_230; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_231; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_232; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_233; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_234; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_235; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_236; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_237; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_238; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_239; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_240; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_241; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_242; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_243; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_244; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_245; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_246; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_247; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_248; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_249; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_250; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_251; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_252; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_253; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_254; // @[AsyncQueue.scala 113:25]
  wire [7:0] _GEN_255; // @[AsyncQueue.scala 113:25]
  wire [7:0] deq_bits_nxt; // @[AsyncQueue.scala 113:25]
  wire  valid_reg_1; // @[AsyncQueue.scala 116:59]
  wire  _T_293; // @[AsyncQueue.scala 117:29]
  wire  _T_298; // @[AsyncQueue.scala 127:37]
  wire  _T_299; // @[AsyncQueue.scala 127:34]
  wire  _T_318; // @[AsyncQueue.scala 139:59]
  wire [7:0] _T_291; // @[ShiftReg.scala 50:24]
  AsyncResetRegVec_w9_i0 ridx_bin ( // @[AsyncResetReg.scala 110:21]
    .clock(ridx_bin_clock),
    .reset(ridx_bin_reset),
    .io_d(ridx_bin_io_d),
    .io_q(ridx_bin_io_q),
    .io_en(ridx_bin_io_en)
  );
  AsyncResetSynchronizerShiftReg_w9_d3_i0 widx_gray ( // @[ShiftReg.scala 47:23]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q)
  );
  SynchronizerShiftReg_w8_d1 deq_bits_reg ( // @[ShiftReg.scala 47:23]
    .clock(deq_bits_reg_clock),
    .io_d(deq_bits_reg_io_d),
    .io_q(deq_bits_reg_io_q)
  );
  AsyncResetRegVec_w1_i0 valid_reg ( // @[AsyncResetReg.scala 110:21]
    .clock(valid_reg_clock),
    .reset(valid_reg_reset),
    .io_d(valid_reg_io_d),
    .io_q(valid_reg_io_q),
    .io_en(valid_reg_io_en)
  );
  AsyncResetRegVec_w9_i0 ridx_gray ( // @[AsyncResetReg.scala 110:21]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q),
    .io_en(ridx_gray_io_en)
  );
  AsyncValidSync_3 AsyncValidSync ( // @[AsyncQueue.scala 124:31]
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_4 AsyncValidSync_1 ( // @[AsyncQueue.scala 125:31]
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_5 AsyncValidSync_2 ( // @[AsyncQueue.scala 126:31]
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  AsyncResetRegVec_w1_i0 AsyncResetRegVec_w1_i0 ( // @[AsyncResetReg.scala 110:21]
    .clock(AsyncResetRegVec_w1_i0_clock),
    .reset(AsyncResetRegVec_w1_i0_reset),
    .io_d(AsyncResetRegVec_w1_i0_io_d),
    .io_q(AsyncResetRegVec_w1_i0_io_q),
    .io_en(AsyncResetRegVec_w1_i0_io_en)
  );
  assign _T_272 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 30:37]
  assign source_ready = AsyncValidSync_2_io_out;
  assign _T_274 = source_ready == 1'h0; // @[AsyncQueue.scala 99:49]
  assign _GEN_256 = {{8'd0}, _T_272}; // @[AsyncQueue.scala 11:47]
  assign _T_279 = ridx_bin_io_q + _GEN_256; // @[AsyncQueue.scala 11:47]
  assign _T_280 = _T_279[8:0]; // @[AsyncQueue.scala 11:47]
  assign _T_281 = _T_274 ? 9'h0 : _T_280; // @[AsyncQueue.scala 11:23]
  assign _T_283 = _T_281 >> 1'h1; // @[AsyncQueue.scala 12:32]
  assign ridx = _T_281 ^ _T_283; // @[AsyncQueue.scala 12:17]
  assign widx = widx_gray_io_q; // @[ShiftReg.scala 50:24]
  assign _T_285 = ridx != widx; // @[AsyncQueue.scala 101:36]
  assign valid = source_ready & _T_285; // @[AsyncQueue.scala 101:28]
  assign _T_286 = ridx[7:0]; // @[AsyncQueue.scala 107:48]
  assign _T_287 = ridx[8]; // @[AsyncQueue.scala 107:67]
  assign _GEN_257 = {{7'd0}, _T_287}; // @[AsyncQueue.scala 107:80]
  assign _T_288 = _GEN_257 << 7; // @[AsyncQueue.scala 107:80]
  assign index = _T_286 ^ _T_288; // @[AsyncQueue.scala 107:60]
  assign _GEN_1 = 8'h1 == index ? io_mem_1 : io_mem_0; // @[AsyncQueue.scala 113:25]
  assign _GEN_2 = 8'h2 == index ? io_mem_2 : _GEN_1; // @[AsyncQueue.scala 113:25]
  assign _GEN_3 = 8'h3 == index ? io_mem_3 : _GEN_2; // @[AsyncQueue.scala 113:25]
  assign _GEN_4 = 8'h4 == index ? io_mem_4 : _GEN_3; // @[AsyncQueue.scala 113:25]
  assign _GEN_5 = 8'h5 == index ? io_mem_5 : _GEN_4; // @[AsyncQueue.scala 113:25]
  assign _GEN_6 = 8'h6 == index ? io_mem_6 : _GEN_5; // @[AsyncQueue.scala 113:25]
  assign _GEN_7 = 8'h7 == index ? io_mem_7 : _GEN_6; // @[AsyncQueue.scala 113:25]
  assign _GEN_8 = 8'h8 == index ? io_mem_8 : _GEN_7; // @[AsyncQueue.scala 113:25]
  assign _GEN_9 = 8'h9 == index ? io_mem_9 : _GEN_8; // @[AsyncQueue.scala 113:25]
  assign _GEN_10 = 8'ha == index ? io_mem_10 : _GEN_9; // @[AsyncQueue.scala 113:25]
  assign _GEN_11 = 8'hb == index ? io_mem_11 : _GEN_10; // @[AsyncQueue.scala 113:25]
  assign _GEN_12 = 8'hc == index ? io_mem_12 : _GEN_11; // @[AsyncQueue.scala 113:25]
  assign _GEN_13 = 8'hd == index ? io_mem_13 : _GEN_12; // @[AsyncQueue.scala 113:25]
  assign _GEN_14 = 8'he == index ? io_mem_14 : _GEN_13; // @[AsyncQueue.scala 113:25]
  assign _GEN_15 = 8'hf == index ? io_mem_15 : _GEN_14; // @[AsyncQueue.scala 113:25]
  assign _GEN_16 = 8'h10 == index ? io_mem_16 : _GEN_15; // @[AsyncQueue.scala 113:25]
  assign _GEN_17 = 8'h11 == index ? io_mem_17 : _GEN_16; // @[AsyncQueue.scala 113:25]
  assign _GEN_18 = 8'h12 == index ? io_mem_18 : _GEN_17; // @[AsyncQueue.scala 113:25]
  assign _GEN_19 = 8'h13 == index ? io_mem_19 : _GEN_18; // @[AsyncQueue.scala 113:25]
  assign _GEN_20 = 8'h14 == index ? io_mem_20 : _GEN_19; // @[AsyncQueue.scala 113:25]
  assign _GEN_21 = 8'h15 == index ? io_mem_21 : _GEN_20; // @[AsyncQueue.scala 113:25]
  assign _GEN_22 = 8'h16 == index ? io_mem_22 : _GEN_21; // @[AsyncQueue.scala 113:25]
  assign _GEN_23 = 8'h17 == index ? io_mem_23 : _GEN_22; // @[AsyncQueue.scala 113:25]
  assign _GEN_24 = 8'h18 == index ? io_mem_24 : _GEN_23; // @[AsyncQueue.scala 113:25]
  assign _GEN_25 = 8'h19 == index ? io_mem_25 : _GEN_24; // @[AsyncQueue.scala 113:25]
  assign _GEN_26 = 8'h1a == index ? io_mem_26 : _GEN_25; // @[AsyncQueue.scala 113:25]
  assign _GEN_27 = 8'h1b == index ? io_mem_27 : _GEN_26; // @[AsyncQueue.scala 113:25]
  assign _GEN_28 = 8'h1c == index ? io_mem_28 : _GEN_27; // @[AsyncQueue.scala 113:25]
  assign _GEN_29 = 8'h1d == index ? io_mem_29 : _GEN_28; // @[AsyncQueue.scala 113:25]
  assign _GEN_30 = 8'h1e == index ? io_mem_30 : _GEN_29; // @[AsyncQueue.scala 113:25]
  assign _GEN_31 = 8'h1f == index ? io_mem_31 : _GEN_30; // @[AsyncQueue.scala 113:25]
  assign _GEN_32 = 8'h20 == index ? io_mem_32 : _GEN_31; // @[AsyncQueue.scala 113:25]
  assign _GEN_33 = 8'h21 == index ? io_mem_33 : _GEN_32; // @[AsyncQueue.scala 113:25]
  assign _GEN_34 = 8'h22 == index ? io_mem_34 : _GEN_33; // @[AsyncQueue.scala 113:25]
  assign _GEN_35 = 8'h23 == index ? io_mem_35 : _GEN_34; // @[AsyncQueue.scala 113:25]
  assign _GEN_36 = 8'h24 == index ? io_mem_36 : _GEN_35; // @[AsyncQueue.scala 113:25]
  assign _GEN_37 = 8'h25 == index ? io_mem_37 : _GEN_36; // @[AsyncQueue.scala 113:25]
  assign _GEN_38 = 8'h26 == index ? io_mem_38 : _GEN_37; // @[AsyncQueue.scala 113:25]
  assign _GEN_39 = 8'h27 == index ? io_mem_39 : _GEN_38; // @[AsyncQueue.scala 113:25]
  assign _GEN_40 = 8'h28 == index ? io_mem_40 : _GEN_39; // @[AsyncQueue.scala 113:25]
  assign _GEN_41 = 8'h29 == index ? io_mem_41 : _GEN_40; // @[AsyncQueue.scala 113:25]
  assign _GEN_42 = 8'h2a == index ? io_mem_42 : _GEN_41; // @[AsyncQueue.scala 113:25]
  assign _GEN_43 = 8'h2b == index ? io_mem_43 : _GEN_42; // @[AsyncQueue.scala 113:25]
  assign _GEN_44 = 8'h2c == index ? io_mem_44 : _GEN_43; // @[AsyncQueue.scala 113:25]
  assign _GEN_45 = 8'h2d == index ? io_mem_45 : _GEN_44; // @[AsyncQueue.scala 113:25]
  assign _GEN_46 = 8'h2e == index ? io_mem_46 : _GEN_45; // @[AsyncQueue.scala 113:25]
  assign _GEN_47 = 8'h2f == index ? io_mem_47 : _GEN_46; // @[AsyncQueue.scala 113:25]
  assign _GEN_48 = 8'h30 == index ? io_mem_48 : _GEN_47; // @[AsyncQueue.scala 113:25]
  assign _GEN_49 = 8'h31 == index ? io_mem_49 : _GEN_48; // @[AsyncQueue.scala 113:25]
  assign _GEN_50 = 8'h32 == index ? io_mem_50 : _GEN_49; // @[AsyncQueue.scala 113:25]
  assign _GEN_51 = 8'h33 == index ? io_mem_51 : _GEN_50; // @[AsyncQueue.scala 113:25]
  assign _GEN_52 = 8'h34 == index ? io_mem_52 : _GEN_51; // @[AsyncQueue.scala 113:25]
  assign _GEN_53 = 8'h35 == index ? io_mem_53 : _GEN_52; // @[AsyncQueue.scala 113:25]
  assign _GEN_54 = 8'h36 == index ? io_mem_54 : _GEN_53; // @[AsyncQueue.scala 113:25]
  assign _GEN_55 = 8'h37 == index ? io_mem_55 : _GEN_54; // @[AsyncQueue.scala 113:25]
  assign _GEN_56 = 8'h38 == index ? io_mem_56 : _GEN_55; // @[AsyncQueue.scala 113:25]
  assign _GEN_57 = 8'h39 == index ? io_mem_57 : _GEN_56; // @[AsyncQueue.scala 113:25]
  assign _GEN_58 = 8'h3a == index ? io_mem_58 : _GEN_57; // @[AsyncQueue.scala 113:25]
  assign _GEN_59 = 8'h3b == index ? io_mem_59 : _GEN_58; // @[AsyncQueue.scala 113:25]
  assign _GEN_60 = 8'h3c == index ? io_mem_60 : _GEN_59; // @[AsyncQueue.scala 113:25]
  assign _GEN_61 = 8'h3d == index ? io_mem_61 : _GEN_60; // @[AsyncQueue.scala 113:25]
  assign _GEN_62 = 8'h3e == index ? io_mem_62 : _GEN_61; // @[AsyncQueue.scala 113:25]
  assign _GEN_63 = 8'h3f == index ? io_mem_63 : _GEN_62; // @[AsyncQueue.scala 113:25]
  assign _GEN_64 = 8'h40 == index ? io_mem_64 : _GEN_63; // @[AsyncQueue.scala 113:25]
  assign _GEN_65 = 8'h41 == index ? io_mem_65 : _GEN_64; // @[AsyncQueue.scala 113:25]
  assign _GEN_66 = 8'h42 == index ? io_mem_66 : _GEN_65; // @[AsyncQueue.scala 113:25]
  assign _GEN_67 = 8'h43 == index ? io_mem_67 : _GEN_66; // @[AsyncQueue.scala 113:25]
  assign _GEN_68 = 8'h44 == index ? io_mem_68 : _GEN_67; // @[AsyncQueue.scala 113:25]
  assign _GEN_69 = 8'h45 == index ? io_mem_69 : _GEN_68; // @[AsyncQueue.scala 113:25]
  assign _GEN_70 = 8'h46 == index ? io_mem_70 : _GEN_69; // @[AsyncQueue.scala 113:25]
  assign _GEN_71 = 8'h47 == index ? io_mem_71 : _GEN_70; // @[AsyncQueue.scala 113:25]
  assign _GEN_72 = 8'h48 == index ? io_mem_72 : _GEN_71; // @[AsyncQueue.scala 113:25]
  assign _GEN_73 = 8'h49 == index ? io_mem_73 : _GEN_72; // @[AsyncQueue.scala 113:25]
  assign _GEN_74 = 8'h4a == index ? io_mem_74 : _GEN_73; // @[AsyncQueue.scala 113:25]
  assign _GEN_75 = 8'h4b == index ? io_mem_75 : _GEN_74; // @[AsyncQueue.scala 113:25]
  assign _GEN_76 = 8'h4c == index ? io_mem_76 : _GEN_75; // @[AsyncQueue.scala 113:25]
  assign _GEN_77 = 8'h4d == index ? io_mem_77 : _GEN_76; // @[AsyncQueue.scala 113:25]
  assign _GEN_78 = 8'h4e == index ? io_mem_78 : _GEN_77; // @[AsyncQueue.scala 113:25]
  assign _GEN_79 = 8'h4f == index ? io_mem_79 : _GEN_78; // @[AsyncQueue.scala 113:25]
  assign _GEN_80 = 8'h50 == index ? io_mem_80 : _GEN_79; // @[AsyncQueue.scala 113:25]
  assign _GEN_81 = 8'h51 == index ? io_mem_81 : _GEN_80; // @[AsyncQueue.scala 113:25]
  assign _GEN_82 = 8'h52 == index ? io_mem_82 : _GEN_81; // @[AsyncQueue.scala 113:25]
  assign _GEN_83 = 8'h53 == index ? io_mem_83 : _GEN_82; // @[AsyncQueue.scala 113:25]
  assign _GEN_84 = 8'h54 == index ? io_mem_84 : _GEN_83; // @[AsyncQueue.scala 113:25]
  assign _GEN_85 = 8'h55 == index ? io_mem_85 : _GEN_84; // @[AsyncQueue.scala 113:25]
  assign _GEN_86 = 8'h56 == index ? io_mem_86 : _GEN_85; // @[AsyncQueue.scala 113:25]
  assign _GEN_87 = 8'h57 == index ? io_mem_87 : _GEN_86; // @[AsyncQueue.scala 113:25]
  assign _GEN_88 = 8'h58 == index ? io_mem_88 : _GEN_87; // @[AsyncQueue.scala 113:25]
  assign _GEN_89 = 8'h59 == index ? io_mem_89 : _GEN_88; // @[AsyncQueue.scala 113:25]
  assign _GEN_90 = 8'h5a == index ? io_mem_90 : _GEN_89; // @[AsyncQueue.scala 113:25]
  assign _GEN_91 = 8'h5b == index ? io_mem_91 : _GEN_90; // @[AsyncQueue.scala 113:25]
  assign _GEN_92 = 8'h5c == index ? io_mem_92 : _GEN_91; // @[AsyncQueue.scala 113:25]
  assign _GEN_93 = 8'h5d == index ? io_mem_93 : _GEN_92; // @[AsyncQueue.scala 113:25]
  assign _GEN_94 = 8'h5e == index ? io_mem_94 : _GEN_93; // @[AsyncQueue.scala 113:25]
  assign _GEN_95 = 8'h5f == index ? io_mem_95 : _GEN_94; // @[AsyncQueue.scala 113:25]
  assign _GEN_96 = 8'h60 == index ? io_mem_96 : _GEN_95; // @[AsyncQueue.scala 113:25]
  assign _GEN_97 = 8'h61 == index ? io_mem_97 : _GEN_96; // @[AsyncQueue.scala 113:25]
  assign _GEN_98 = 8'h62 == index ? io_mem_98 : _GEN_97; // @[AsyncQueue.scala 113:25]
  assign _GEN_99 = 8'h63 == index ? io_mem_99 : _GEN_98; // @[AsyncQueue.scala 113:25]
  assign _GEN_100 = 8'h64 == index ? io_mem_100 : _GEN_99; // @[AsyncQueue.scala 113:25]
  assign _GEN_101 = 8'h65 == index ? io_mem_101 : _GEN_100; // @[AsyncQueue.scala 113:25]
  assign _GEN_102 = 8'h66 == index ? io_mem_102 : _GEN_101; // @[AsyncQueue.scala 113:25]
  assign _GEN_103 = 8'h67 == index ? io_mem_103 : _GEN_102; // @[AsyncQueue.scala 113:25]
  assign _GEN_104 = 8'h68 == index ? io_mem_104 : _GEN_103; // @[AsyncQueue.scala 113:25]
  assign _GEN_105 = 8'h69 == index ? io_mem_105 : _GEN_104; // @[AsyncQueue.scala 113:25]
  assign _GEN_106 = 8'h6a == index ? io_mem_106 : _GEN_105; // @[AsyncQueue.scala 113:25]
  assign _GEN_107 = 8'h6b == index ? io_mem_107 : _GEN_106; // @[AsyncQueue.scala 113:25]
  assign _GEN_108 = 8'h6c == index ? io_mem_108 : _GEN_107; // @[AsyncQueue.scala 113:25]
  assign _GEN_109 = 8'h6d == index ? io_mem_109 : _GEN_108; // @[AsyncQueue.scala 113:25]
  assign _GEN_110 = 8'h6e == index ? io_mem_110 : _GEN_109; // @[AsyncQueue.scala 113:25]
  assign _GEN_111 = 8'h6f == index ? io_mem_111 : _GEN_110; // @[AsyncQueue.scala 113:25]
  assign _GEN_112 = 8'h70 == index ? io_mem_112 : _GEN_111; // @[AsyncQueue.scala 113:25]
  assign _GEN_113 = 8'h71 == index ? io_mem_113 : _GEN_112; // @[AsyncQueue.scala 113:25]
  assign _GEN_114 = 8'h72 == index ? io_mem_114 : _GEN_113; // @[AsyncQueue.scala 113:25]
  assign _GEN_115 = 8'h73 == index ? io_mem_115 : _GEN_114; // @[AsyncQueue.scala 113:25]
  assign _GEN_116 = 8'h74 == index ? io_mem_116 : _GEN_115; // @[AsyncQueue.scala 113:25]
  assign _GEN_117 = 8'h75 == index ? io_mem_117 : _GEN_116; // @[AsyncQueue.scala 113:25]
  assign _GEN_118 = 8'h76 == index ? io_mem_118 : _GEN_117; // @[AsyncQueue.scala 113:25]
  assign _GEN_119 = 8'h77 == index ? io_mem_119 : _GEN_118; // @[AsyncQueue.scala 113:25]
  assign _GEN_120 = 8'h78 == index ? io_mem_120 : _GEN_119; // @[AsyncQueue.scala 113:25]
  assign _GEN_121 = 8'h79 == index ? io_mem_121 : _GEN_120; // @[AsyncQueue.scala 113:25]
  assign _GEN_122 = 8'h7a == index ? io_mem_122 : _GEN_121; // @[AsyncQueue.scala 113:25]
  assign _GEN_123 = 8'h7b == index ? io_mem_123 : _GEN_122; // @[AsyncQueue.scala 113:25]
  assign _GEN_124 = 8'h7c == index ? io_mem_124 : _GEN_123; // @[AsyncQueue.scala 113:25]
  assign _GEN_125 = 8'h7d == index ? io_mem_125 : _GEN_124; // @[AsyncQueue.scala 113:25]
  assign _GEN_126 = 8'h7e == index ? io_mem_126 : _GEN_125; // @[AsyncQueue.scala 113:25]
  assign _GEN_127 = 8'h7f == index ? io_mem_127 : _GEN_126; // @[AsyncQueue.scala 113:25]
  assign _GEN_128 = 8'h80 == index ? io_mem_128 : _GEN_127; // @[AsyncQueue.scala 113:25]
  assign _GEN_129 = 8'h81 == index ? io_mem_129 : _GEN_128; // @[AsyncQueue.scala 113:25]
  assign _GEN_130 = 8'h82 == index ? io_mem_130 : _GEN_129; // @[AsyncQueue.scala 113:25]
  assign _GEN_131 = 8'h83 == index ? io_mem_131 : _GEN_130; // @[AsyncQueue.scala 113:25]
  assign _GEN_132 = 8'h84 == index ? io_mem_132 : _GEN_131; // @[AsyncQueue.scala 113:25]
  assign _GEN_133 = 8'h85 == index ? io_mem_133 : _GEN_132; // @[AsyncQueue.scala 113:25]
  assign _GEN_134 = 8'h86 == index ? io_mem_134 : _GEN_133; // @[AsyncQueue.scala 113:25]
  assign _GEN_135 = 8'h87 == index ? io_mem_135 : _GEN_134; // @[AsyncQueue.scala 113:25]
  assign _GEN_136 = 8'h88 == index ? io_mem_136 : _GEN_135; // @[AsyncQueue.scala 113:25]
  assign _GEN_137 = 8'h89 == index ? io_mem_137 : _GEN_136; // @[AsyncQueue.scala 113:25]
  assign _GEN_138 = 8'h8a == index ? io_mem_138 : _GEN_137; // @[AsyncQueue.scala 113:25]
  assign _GEN_139 = 8'h8b == index ? io_mem_139 : _GEN_138; // @[AsyncQueue.scala 113:25]
  assign _GEN_140 = 8'h8c == index ? io_mem_140 : _GEN_139; // @[AsyncQueue.scala 113:25]
  assign _GEN_141 = 8'h8d == index ? io_mem_141 : _GEN_140; // @[AsyncQueue.scala 113:25]
  assign _GEN_142 = 8'h8e == index ? io_mem_142 : _GEN_141; // @[AsyncQueue.scala 113:25]
  assign _GEN_143 = 8'h8f == index ? io_mem_143 : _GEN_142; // @[AsyncQueue.scala 113:25]
  assign _GEN_144 = 8'h90 == index ? io_mem_144 : _GEN_143; // @[AsyncQueue.scala 113:25]
  assign _GEN_145 = 8'h91 == index ? io_mem_145 : _GEN_144; // @[AsyncQueue.scala 113:25]
  assign _GEN_146 = 8'h92 == index ? io_mem_146 : _GEN_145; // @[AsyncQueue.scala 113:25]
  assign _GEN_147 = 8'h93 == index ? io_mem_147 : _GEN_146; // @[AsyncQueue.scala 113:25]
  assign _GEN_148 = 8'h94 == index ? io_mem_148 : _GEN_147; // @[AsyncQueue.scala 113:25]
  assign _GEN_149 = 8'h95 == index ? io_mem_149 : _GEN_148; // @[AsyncQueue.scala 113:25]
  assign _GEN_150 = 8'h96 == index ? io_mem_150 : _GEN_149; // @[AsyncQueue.scala 113:25]
  assign _GEN_151 = 8'h97 == index ? io_mem_151 : _GEN_150; // @[AsyncQueue.scala 113:25]
  assign _GEN_152 = 8'h98 == index ? io_mem_152 : _GEN_151; // @[AsyncQueue.scala 113:25]
  assign _GEN_153 = 8'h99 == index ? io_mem_153 : _GEN_152; // @[AsyncQueue.scala 113:25]
  assign _GEN_154 = 8'h9a == index ? io_mem_154 : _GEN_153; // @[AsyncQueue.scala 113:25]
  assign _GEN_155 = 8'h9b == index ? io_mem_155 : _GEN_154; // @[AsyncQueue.scala 113:25]
  assign _GEN_156 = 8'h9c == index ? io_mem_156 : _GEN_155; // @[AsyncQueue.scala 113:25]
  assign _GEN_157 = 8'h9d == index ? io_mem_157 : _GEN_156; // @[AsyncQueue.scala 113:25]
  assign _GEN_158 = 8'h9e == index ? io_mem_158 : _GEN_157; // @[AsyncQueue.scala 113:25]
  assign _GEN_159 = 8'h9f == index ? io_mem_159 : _GEN_158; // @[AsyncQueue.scala 113:25]
  assign _GEN_160 = 8'ha0 == index ? io_mem_160 : _GEN_159; // @[AsyncQueue.scala 113:25]
  assign _GEN_161 = 8'ha1 == index ? io_mem_161 : _GEN_160; // @[AsyncQueue.scala 113:25]
  assign _GEN_162 = 8'ha2 == index ? io_mem_162 : _GEN_161; // @[AsyncQueue.scala 113:25]
  assign _GEN_163 = 8'ha3 == index ? io_mem_163 : _GEN_162; // @[AsyncQueue.scala 113:25]
  assign _GEN_164 = 8'ha4 == index ? io_mem_164 : _GEN_163; // @[AsyncQueue.scala 113:25]
  assign _GEN_165 = 8'ha5 == index ? io_mem_165 : _GEN_164; // @[AsyncQueue.scala 113:25]
  assign _GEN_166 = 8'ha6 == index ? io_mem_166 : _GEN_165; // @[AsyncQueue.scala 113:25]
  assign _GEN_167 = 8'ha7 == index ? io_mem_167 : _GEN_166; // @[AsyncQueue.scala 113:25]
  assign _GEN_168 = 8'ha8 == index ? io_mem_168 : _GEN_167; // @[AsyncQueue.scala 113:25]
  assign _GEN_169 = 8'ha9 == index ? io_mem_169 : _GEN_168; // @[AsyncQueue.scala 113:25]
  assign _GEN_170 = 8'haa == index ? io_mem_170 : _GEN_169; // @[AsyncQueue.scala 113:25]
  assign _GEN_171 = 8'hab == index ? io_mem_171 : _GEN_170; // @[AsyncQueue.scala 113:25]
  assign _GEN_172 = 8'hac == index ? io_mem_172 : _GEN_171; // @[AsyncQueue.scala 113:25]
  assign _GEN_173 = 8'had == index ? io_mem_173 : _GEN_172; // @[AsyncQueue.scala 113:25]
  assign _GEN_174 = 8'hae == index ? io_mem_174 : _GEN_173; // @[AsyncQueue.scala 113:25]
  assign _GEN_175 = 8'haf == index ? io_mem_175 : _GEN_174; // @[AsyncQueue.scala 113:25]
  assign _GEN_176 = 8'hb0 == index ? io_mem_176 : _GEN_175; // @[AsyncQueue.scala 113:25]
  assign _GEN_177 = 8'hb1 == index ? io_mem_177 : _GEN_176; // @[AsyncQueue.scala 113:25]
  assign _GEN_178 = 8'hb2 == index ? io_mem_178 : _GEN_177; // @[AsyncQueue.scala 113:25]
  assign _GEN_179 = 8'hb3 == index ? io_mem_179 : _GEN_178; // @[AsyncQueue.scala 113:25]
  assign _GEN_180 = 8'hb4 == index ? io_mem_180 : _GEN_179; // @[AsyncQueue.scala 113:25]
  assign _GEN_181 = 8'hb5 == index ? io_mem_181 : _GEN_180; // @[AsyncQueue.scala 113:25]
  assign _GEN_182 = 8'hb6 == index ? io_mem_182 : _GEN_181; // @[AsyncQueue.scala 113:25]
  assign _GEN_183 = 8'hb7 == index ? io_mem_183 : _GEN_182; // @[AsyncQueue.scala 113:25]
  assign _GEN_184 = 8'hb8 == index ? io_mem_184 : _GEN_183; // @[AsyncQueue.scala 113:25]
  assign _GEN_185 = 8'hb9 == index ? io_mem_185 : _GEN_184; // @[AsyncQueue.scala 113:25]
  assign _GEN_186 = 8'hba == index ? io_mem_186 : _GEN_185; // @[AsyncQueue.scala 113:25]
  assign _GEN_187 = 8'hbb == index ? io_mem_187 : _GEN_186; // @[AsyncQueue.scala 113:25]
  assign _GEN_188 = 8'hbc == index ? io_mem_188 : _GEN_187; // @[AsyncQueue.scala 113:25]
  assign _GEN_189 = 8'hbd == index ? io_mem_189 : _GEN_188; // @[AsyncQueue.scala 113:25]
  assign _GEN_190 = 8'hbe == index ? io_mem_190 : _GEN_189; // @[AsyncQueue.scala 113:25]
  assign _GEN_191 = 8'hbf == index ? io_mem_191 : _GEN_190; // @[AsyncQueue.scala 113:25]
  assign _GEN_192 = 8'hc0 == index ? io_mem_192 : _GEN_191; // @[AsyncQueue.scala 113:25]
  assign _GEN_193 = 8'hc1 == index ? io_mem_193 : _GEN_192; // @[AsyncQueue.scala 113:25]
  assign _GEN_194 = 8'hc2 == index ? io_mem_194 : _GEN_193; // @[AsyncQueue.scala 113:25]
  assign _GEN_195 = 8'hc3 == index ? io_mem_195 : _GEN_194; // @[AsyncQueue.scala 113:25]
  assign _GEN_196 = 8'hc4 == index ? io_mem_196 : _GEN_195; // @[AsyncQueue.scala 113:25]
  assign _GEN_197 = 8'hc5 == index ? io_mem_197 : _GEN_196; // @[AsyncQueue.scala 113:25]
  assign _GEN_198 = 8'hc6 == index ? io_mem_198 : _GEN_197; // @[AsyncQueue.scala 113:25]
  assign _GEN_199 = 8'hc7 == index ? io_mem_199 : _GEN_198; // @[AsyncQueue.scala 113:25]
  assign _GEN_200 = 8'hc8 == index ? io_mem_200 : _GEN_199; // @[AsyncQueue.scala 113:25]
  assign _GEN_201 = 8'hc9 == index ? io_mem_201 : _GEN_200; // @[AsyncQueue.scala 113:25]
  assign _GEN_202 = 8'hca == index ? io_mem_202 : _GEN_201; // @[AsyncQueue.scala 113:25]
  assign _GEN_203 = 8'hcb == index ? io_mem_203 : _GEN_202; // @[AsyncQueue.scala 113:25]
  assign _GEN_204 = 8'hcc == index ? io_mem_204 : _GEN_203; // @[AsyncQueue.scala 113:25]
  assign _GEN_205 = 8'hcd == index ? io_mem_205 : _GEN_204; // @[AsyncQueue.scala 113:25]
  assign _GEN_206 = 8'hce == index ? io_mem_206 : _GEN_205; // @[AsyncQueue.scala 113:25]
  assign _GEN_207 = 8'hcf == index ? io_mem_207 : _GEN_206; // @[AsyncQueue.scala 113:25]
  assign _GEN_208 = 8'hd0 == index ? io_mem_208 : _GEN_207; // @[AsyncQueue.scala 113:25]
  assign _GEN_209 = 8'hd1 == index ? io_mem_209 : _GEN_208; // @[AsyncQueue.scala 113:25]
  assign _GEN_210 = 8'hd2 == index ? io_mem_210 : _GEN_209; // @[AsyncQueue.scala 113:25]
  assign _GEN_211 = 8'hd3 == index ? io_mem_211 : _GEN_210; // @[AsyncQueue.scala 113:25]
  assign _GEN_212 = 8'hd4 == index ? io_mem_212 : _GEN_211; // @[AsyncQueue.scala 113:25]
  assign _GEN_213 = 8'hd5 == index ? io_mem_213 : _GEN_212; // @[AsyncQueue.scala 113:25]
  assign _GEN_214 = 8'hd6 == index ? io_mem_214 : _GEN_213; // @[AsyncQueue.scala 113:25]
  assign _GEN_215 = 8'hd7 == index ? io_mem_215 : _GEN_214; // @[AsyncQueue.scala 113:25]
  assign _GEN_216 = 8'hd8 == index ? io_mem_216 : _GEN_215; // @[AsyncQueue.scala 113:25]
  assign _GEN_217 = 8'hd9 == index ? io_mem_217 : _GEN_216; // @[AsyncQueue.scala 113:25]
  assign _GEN_218 = 8'hda == index ? io_mem_218 : _GEN_217; // @[AsyncQueue.scala 113:25]
  assign _GEN_219 = 8'hdb == index ? io_mem_219 : _GEN_218; // @[AsyncQueue.scala 113:25]
  assign _GEN_220 = 8'hdc == index ? io_mem_220 : _GEN_219; // @[AsyncQueue.scala 113:25]
  assign _GEN_221 = 8'hdd == index ? io_mem_221 : _GEN_220; // @[AsyncQueue.scala 113:25]
  assign _GEN_222 = 8'hde == index ? io_mem_222 : _GEN_221; // @[AsyncQueue.scala 113:25]
  assign _GEN_223 = 8'hdf == index ? io_mem_223 : _GEN_222; // @[AsyncQueue.scala 113:25]
  assign _GEN_224 = 8'he0 == index ? io_mem_224 : _GEN_223; // @[AsyncQueue.scala 113:25]
  assign _GEN_225 = 8'he1 == index ? io_mem_225 : _GEN_224; // @[AsyncQueue.scala 113:25]
  assign _GEN_226 = 8'he2 == index ? io_mem_226 : _GEN_225; // @[AsyncQueue.scala 113:25]
  assign _GEN_227 = 8'he3 == index ? io_mem_227 : _GEN_226; // @[AsyncQueue.scala 113:25]
  assign _GEN_228 = 8'he4 == index ? io_mem_228 : _GEN_227; // @[AsyncQueue.scala 113:25]
  assign _GEN_229 = 8'he5 == index ? io_mem_229 : _GEN_228; // @[AsyncQueue.scala 113:25]
  assign _GEN_230 = 8'he6 == index ? io_mem_230 : _GEN_229; // @[AsyncQueue.scala 113:25]
  assign _GEN_231 = 8'he7 == index ? io_mem_231 : _GEN_230; // @[AsyncQueue.scala 113:25]
  assign _GEN_232 = 8'he8 == index ? io_mem_232 : _GEN_231; // @[AsyncQueue.scala 113:25]
  assign _GEN_233 = 8'he9 == index ? io_mem_233 : _GEN_232; // @[AsyncQueue.scala 113:25]
  assign _GEN_234 = 8'hea == index ? io_mem_234 : _GEN_233; // @[AsyncQueue.scala 113:25]
  assign _GEN_235 = 8'heb == index ? io_mem_235 : _GEN_234; // @[AsyncQueue.scala 113:25]
  assign _GEN_236 = 8'hec == index ? io_mem_236 : _GEN_235; // @[AsyncQueue.scala 113:25]
  assign _GEN_237 = 8'hed == index ? io_mem_237 : _GEN_236; // @[AsyncQueue.scala 113:25]
  assign _GEN_238 = 8'hee == index ? io_mem_238 : _GEN_237; // @[AsyncQueue.scala 113:25]
  assign _GEN_239 = 8'hef == index ? io_mem_239 : _GEN_238; // @[AsyncQueue.scala 113:25]
  assign _GEN_240 = 8'hf0 == index ? io_mem_240 : _GEN_239; // @[AsyncQueue.scala 113:25]
  assign _GEN_241 = 8'hf1 == index ? io_mem_241 : _GEN_240; // @[AsyncQueue.scala 113:25]
  assign _GEN_242 = 8'hf2 == index ? io_mem_242 : _GEN_241; // @[AsyncQueue.scala 113:25]
  assign _GEN_243 = 8'hf3 == index ? io_mem_243 : _GEN_242; // @[AsyncQueue.scala 113:25]
  assign _GEN_244 = 8'hf4 == index ? io_mem_244 : _GEN_243; // @[AsyncQueue.scala 113:25]
  assign _GEN_245 = 8'hf5 == index ? io_mem_245 : _GEN_244; // @[AsyncQueue.scala 113:25]
  assign _GEN_246 = 8'hf6 == index ? io_mem_246 : _GEN_245; // @[AsyncQueue.scala 113:25]
  assign _GEN_247 = 8'hf7 == index ? io_mem_247 : _GEN_246; // @[AsyncQueue.scala 113:25]
  assign _GEN_248 = 8'hf8 == index ? io_mem_248 : _GEN_247; // @[AsyncQueue.scala 113:25]
  assign _GEN_249 = 8'hf9 == index ? io_mem_249 : _GEN_248; // @[AsyncQueue.scala 113:25]
  assign _GEN_250 = 8'hfa == index ? io_mem_250 : _GEN_249; // @[AsyncQueue.scala 113:25]
  assign _GEN_251 = 8'hfb == index ? io_mem_251 : _GEN_250; // @[AsyncQueue.scala 113:25]
  assign _GEN_252 = 8'hfc == index ? io_mem_252 : _GEN_251; // @[AsyncQueue.scala 113:25]
  assign _GEN_253 = 8'hfd == index ? io_mem_253 : _GEN_252; // @[AsyncQueue.scala 113:25]
  assign _GEN_254 = 8'hfe == index ? io_mem_254 : _GEN_253; // @[AsyncQueue.scala 113:25]
  assign _GEN_255 = 8'hff == index ? io_mem_255 : _GEN_254; // @[AsyncQueue.scala 113:25]
  assign deq_bits_nxt = valid ? _GEN_255 : io_deq_bits; // @[AsyncQueue.scala 113:25]
  assign valid_reg_1 = valid_reg_io_q; // @[AsyncQueue.scala 116:59]
  assign _T_293 = valid_reg_1 & source_ready; // @[AsyncQueue.scala 117:29]
  assign _T_298 = io_source_reset_n == 1'h0; // @[AsyncQueue.scala 127:37]
  assign _T_299 = reset | _T_298; // @[AsyncQueue.scala 127:34]
  assign _T_318 = io_widx == io_ridx; // @[AsyncQueue.scala 139:59]
  assign _T_291 = deq_bits_reg_io_q; // @[ShiftReg.scala 50:24]
  assign io_deq_valid = _T_293;
  assign io_deq_bits = _T_291;
  assign io_ridx = ridx_gray_io_q;
  assign io_ridx_valid = AsyncValidSync_io_out;
  assign ridx_bin_clock = clock;
  assign ridx_bin_reset = reset;
  assign ridx_bin_io_d = _T_281;
  assign ridx_bin_io_en = 1'h1;
  assign widx_gray_clock = clock;
  assign widx_gray_reset = reset;
  assign widx_gray_io_d = io_widx;
  assign deq_bits_reg_clock = clock;
  assign deq_bits_reg_io_d = deq_bits_nxt;
  assign valid_reg_clock = clock;
  assign valid_reg_reset = reset;
  assign valid_reg_io_d = valid;
  assign valid_reg_io_en = 1'h1;
  assign ridx_gray_clock = clock;
  assign ridx_gray_reset = reset;
  assign ridx_gray_io_d = ridx;
  assign ridx_gray_io_en = 1'h1;
  assign AsyncValidSync_clock = clock;
  assign AsyncValidSync_reset = _T_299;
  assign AsyncValidSync_1_clock = clock;
  assign AsyncValidSync_1_reset = _T_299;
  assign AsyncValidSync_1_io_in = io_widx_valid;
  assign AsyncValidSync_2_clock = clock;
  assign AsyncValidSync_2_reset = reset;
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out;
  assign AsyncResetRegVec_w1_i0_clock = clock;
  assign AsyncResetRegVec_w1_i0_reset = reset;
  assign AsyncResetRegVec_w1_i0_io_d = _T_318;
  assign AsyncResetRegVec_w1_i0_io_en = 1'h1;
endmodule
module AsyncQueue_1(
  input        io_enq_clock,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_clock,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits
);
  wire  source_clock; // @[AsyncQueue.scala 155:22]
  wire  source_reset; // @[AsyncQueue.scala 155:22]
  wire  source_io_enq_ready; // @[AsyncQueue.scala 155:22]
  wire  source_io_enq_valid; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_enq_bits; // @[AsyncQueue.scala 155:22]
  wire [8:0] source_io_ridx; // @[AsyncQueue.scala 155:22]
  wire [8:0] source_io_widx; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_0; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_1; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_2; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_3; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_4; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_5; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_6; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_7; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_8; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_9; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_10; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_11; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_12; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_13; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_14; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_15; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_16; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_17; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_18; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_19; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_20; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_21; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_22; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_23; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_24; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_25; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_26; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_27; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_28; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_29; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_30; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_31; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_32; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_33; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_34; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_35; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_36; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_37; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_38; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_39; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_40; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_41; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_42; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_43; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_44; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_45; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_46; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_47; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_48; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_49; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_50; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_51; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_52; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_53; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_54; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_55; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_56; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_57; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_58; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_59; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_60; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_61; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_62; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_63; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_64; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_65; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_66; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_67; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_68; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_69; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_70; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_71; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_72; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_73; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_74; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_75; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_76; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_77; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_78; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_79; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_80; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_81; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_82; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_83; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_84; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_85; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_86; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_87; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_88; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_89; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_90; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_91; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_92; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_93; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_94; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_95; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_96; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_97; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_98; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_99; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_100; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_101; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_102; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_103; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_104; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_105; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_106; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_107; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_108; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_109; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_110; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_111; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_112; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_113; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_114; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_115; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_116; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_117; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_118; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_119; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_120; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_121; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_122; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_123; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_124; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_125; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_126; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_127; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_128; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_129; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_130; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_131; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_132; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_133; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_134; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_135; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_136; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_137; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_138; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_139; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_140; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_141; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_142; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_143; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_144; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_145; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_146; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_147; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_148; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_149; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_150; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_151; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_152; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_153; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_154; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_155; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_156; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_157; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_158; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_159; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_160; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_161; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_162; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_163; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_164; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_165; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_166; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_167; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_168; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_169; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_170; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_171; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_172; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_173; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_174; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_175; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_176; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_177; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_178; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_179; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_180; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_181; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_182; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_183; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_184; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_185; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_186; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_187; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_188; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_189; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_190; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_191; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_192; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_193; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_194; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_195; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_196; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_197; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_198; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_199; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_200; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_201; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_202; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_203; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_204; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_205; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_206; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_207; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_208; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_209; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_210; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_211; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_212; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_213; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_214; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_215; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_216; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_217; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_218; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_219; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_220; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_221; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_222; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_223; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_224; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_225; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_226; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_227; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_228; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_229; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_230; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_231; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_232; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_233; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_234; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_235; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_236; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_237; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_238; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_239; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_240; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_241; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_242; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_243; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_244; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_245; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_246; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_247; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_248; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_249; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_250; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_251; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_252; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_253; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_254; // @[AsyncQueue.scala 155:22]
  wire [7:0] source_io_mem_255; // @[AsyncQueue.scala 155:22]
  wire  source_io_sink_reset_n; // @[AsyncQueue.scala 155:22]
  wire  source_io_ridx_valid; // @[AsyncQueue.scala 155:22]
  wire  source_io_widx_valid; // @[AsyncQueue.scala 155:22]
  wire  sink_clock; // @[AsyncQueue.scala 156:22]
  wire  sink_reset; // @[AsyncQueue.scala 156:22]
  wire  sink_io_deq_ready; // @[AsyncQueue.scala 156:22]
  wire  sink_io_deq_valid; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_deq_bits; // @[AsyncQueue.scala 156:22]
  wire [8:0] sink_io_ridx; // @[AsyncQueue.scala 156:22]
  wire [8:0] sink_io_widx; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_0; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_1; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_2; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_3; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_4; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_5; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_6; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_7; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_8; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_9; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_10; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_11; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_12; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_13; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_14; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_15; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_16; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_17; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_18; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_19; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_20; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_21; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_22; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_23; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_24; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_25; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_26; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_27; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_28; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_29; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_30; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_31; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_32; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_33; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_34; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_35; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_36; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_37; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_38; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_39; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_40; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_41; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_42; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_43; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_44; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_45; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_46; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_47; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_48; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_49; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_50; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_51; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_52; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_53; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_54; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_55; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_56; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_57; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_58; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_59; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_60; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_61; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_62; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_63; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_64; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_65; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_66; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_67; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_68; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_69; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_70; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_71; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_72; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_73; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_74; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_75; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_76; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_77; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_78; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_79; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_80; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_81; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_82; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_83; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_84; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_85; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_86; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_87; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_88; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_89; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_90; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_91; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_92; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_93; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_94; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_95; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_96; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_97; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_98; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_99; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_100; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_101; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_102; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_103; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_104; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_105; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_106; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_107; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_108; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_109; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_110; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_111; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_112; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_113; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_114; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_115; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_116; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_117; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_118; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_119; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_120; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_121; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_122; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_123; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_124; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_125; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_126; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_127; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_128; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_129; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_130; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_131; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_132; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_133; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_134; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_135; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_136; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_137; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_138; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_139; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_140; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_141; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_142; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_143; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_144; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_145; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_146; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_147; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_148; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_149; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_150; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_151; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_152; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_153; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_154; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_155; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_156; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_157; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_158; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_159; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_160; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_161; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_162; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_163; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_164; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_165; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_166; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_167; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_168; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_169; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_170; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_171; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_172; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_173; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_174; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_175; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_176; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_177; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_178; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_179; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_180; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_181; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_182; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_183; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_184; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_185; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_186; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_187; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_188; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_189; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_190; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_191; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_192; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_193; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_194; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_195; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_196; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_197; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_198; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_199; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_200; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_201; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_202; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_203; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_204; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_205; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_206; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_207; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_208; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_209; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_210; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_211; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_212; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_213; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_214; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_215; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_216; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_217; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_218; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_219; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_220; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_221; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_222; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_223; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_224; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_225; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_226; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_227; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_228; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_229; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_230; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_231; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_232; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_233; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_234; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_235; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_236; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_237; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_238; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_239; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_240; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_241; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_242; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_243; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_244; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_245; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_246; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_247; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_248; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_249; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_250; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_251; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_252; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_253; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_254; // @[AsyncQueue.scala 156:22]
  wire [7:0] sink_io_mem_255; // @[AsyncQueue.scala 156:22]
  wire  sink_io_source_reset_n; // @[AsyncQueue.scala 156:22]
  wire  sink_io_ridx_valid; // @[AsyncQueue.scala 156:22]
  wire  sink_io_widx_valid; // @[AsyncQueue.scala 156:22]
  AsyncQueueSource_1 source ( // @[AsyncQueue.scala 155:22]
    .clock(source_clock),
    .reset(source_reset),
    .io_enq_ready(source_io_enq_ready),
    .io_enq_valid(source_io_enq_valid),
    .io_enq_bits(source_io_enq_bits),
    .io_ridx(source_io_ridx),
    .io_widx(source_io_widx),
    .io_mem_0(source_io_mem_0),
    .io_mem_1(source_io_mem_1),
    .io_mem_2(source_io_mem_2),
    .io_mem_3(source_io_mem_3),
    .io_mem_4(source_io_mem_4),
    .io_mem_5(source_io_mem_5),
    .io_mem_6(source_io_mem_6),
    .io_mem_7(source_io_mem_7),
    .io_mem_8(source_io_mem_8),
    .io_mem_9(source_io_mem_9),
    .io_mem_10(source_io_mem_10),
    .io_mem_11(source_io_mem_11),
    .io_mem_12(source_io_mem_12),
    .io_mem_13(source_io_mem_13),
    .io_mem_14(source_io_mem_14),
    .io_mem_15(source_io_mem_15),
    .io_mem_16(source_io_mem_16),
    .io_mem_17(source_io_mem_17),
    .io_mem_18(source_io_mem_18),
    .io_mem_19(source_io_mem_19),
    .io_mem_20(source_io_mem_20),
    .io_mem_21(source_io_mem_21),
    .io_mem_22(source_io_mem_22),
    .io_mem_23(source_io_mem_23),
    .io_mem_24(source_io_mem_24),
    .io_mem_25(source_io_mem_25),
    .io_mem_26(source_io_mem_26),
    .io_mem_27(source_io_mem_27),
    .io_mem_28(source_io_mem_28),
    .io_mem_29(source_io_mem_29),
    .io_mem_30(source_io_mem_30),
    .io_mem_31(source_io_mem_31),
    .io_mem_32(source_io_mem_32),
    .io_mem_33(source_io_mem_33),
    .io_mem_34(source_io_mem_34),
    .io_mem_35(source_io_mem_35),
    .io_mem_36(source_io_mem_36),
    .io_mem_37(source_io_mem_37),
    .io_mem_38(source_io_mem_38),
    .io_mem_39(source_io_mem_39),
    .io_mem_40(source_io_mem_40),
    .io_mem_41(source_io_mem_41),
    .io_mem_42(source_io_mem_42),
    .io_mem_43(source_io_mem_43),
    .io_mem_44(source_io_mem_44),
    .io_mem_45(source_io_mem_45),
    .io_mem_46(source_io_mem_46),
    .io_mem_47(source_io_mem_47),
    .io_mem_48(source_io_mem_48),
    .io_mem_49(source_io_mem_49),
    .io_mem_50(source_io_mem_50),
    .io_mem_51(source_io_mem_51),
    .io_mem_52(source_io_mem_52),
    .io_mem_53(source_io_mem_53),
    .io_mem_54(source_io_mem_54),
    .io_mem_55(source_io_mem_55),
    .io_mem_56(source_io_mem_56),
    .io_mem_57(source_io_mem_57),
    .io_mem_58(source_io_mem_58),
    .io_mem_59(source_io_mem_59),
    .io_mem_60(source_io_mem_60),
    .io_mem_61(source_io_mem_61),
    .io_mem_62(source_io_mem_62),
    .io_mem_63(source_io_mem_63),
    .io_mem_64(source_io_mem_64),
    .io_mem_65(source_io_mem_65),
    .io_mem_66(source_io_mem_66),
    .io_mem_67(source_io_mem_67),
    .io_mem_68(source_io_mem_68),
    .io_mem_69(source_io_mem_69),
    .io_mem_70(source_io_mem_70),
    .io_mem_71(source_io_mem_71),
    .io_mem_72(source_io_mem_72),
    .io_mem_73(source_io_mem_73),
    .io_mem_74(source_io_mem_74),
    .io_mem_75(source_io_mem_75),
    .io_mem_76(source_io_mem_76),
    .io_mem_77(source_io_mem_77),
    .io_mem_78(source_io_mem_78),
    .io_mem_79(source_io_mem_79),
    .io_mem_80(source_io_mem_80),
    .io_mem_81(source_io_mem_81),
    .io_mem_82(source_io_mem_82),
    .io_mem_83(source_io_mem_83),
    .io_mem_84(source_io_mem_84),
    .io_mem_85(source_io_mem_85),
    .io_mem_86(source_io_mem_86),
    .io_mem_87(source_io_mem_87),
    .io_mem_88(source_io_mem_88),
    .io_mem_89(source_io_mem_89),
    .io_mem_90(source_io_mem_90),
    .io_mem_91(source_io_mem_91),
    .io_mem_92(source_io_mem_92),
    .io_mem_93(source_io_mem_93),
    .io_mem_94(source_io_mem_94),
    .io_mem_95(source_io_mem_95),
    .io_mem_96(source_io_mem_96),
    .io_mem_97(source_io_mem_97),
    .io_mem_98(source_io_mem_98),
    .io_mem_99(source_io_mem_99),
    .io_mem_100(source_io_mem_100),
    .io_mem_101(source_io_mem_101),
    .io_mem_102(source_io_mem_102),
    .io_mem_103(source_io_mem_103),
    .io_mem_104(source_io_mem_104),
    .io_mem_105(source_io_mem_105),
    .io_mem_106(source_io_mem_106),
    .io_mem_107(source_io_mem_107),
    .io_mem_108(source_io_mem_108),
    .io_mem_109(source_io_mem_109),
    .io_mem_110(source_io_mem_110),
    .io_mem_111(source_io_mem_111),
    .io_mem_112(source_io_mem_112),
    .io_mem_113(source_io_mem_113),
    .io_mem_114(source_io_mem_114),
    .io_mem_115(source_io_mem_115),
    .io_mem_116(source_io_mem_116),
    .io_mem_117(source_io_mem_117),
    .io_mem_118(source_io_mem_118),
    .io_mem_119(source_io_mem_119),
    .io_mem_120(source_io_mem_120),
    .io_mem_121(source_io_mem_121),
    .io_mem_122(source_io_mem_122),
    .io_mem_123(source_io_mem_123),
    .io_mem_124(source_io_mem_124),
    .io_mem_125(source_io_mem_125),
    .io_mem_126(source_io_mem_126),
    .io_mem_127(source_io_mem_127),
    .io_mem_128(source_io_mem_128),
    .io_mem_129(source_io_mem_129),
    .io_mem_130(source_io_mem_130),
    .io_mem_131(source_io_mem_131),
    .io_mem_132(source_io_mem_132),
    .io_mem_133(source_io_mem_133),
    .io_mem_134(source_io_mem_134),
    .io_mem_135(source_io_mem_135),
    .io_mem_136(source_io_mem_136),
    .io_mem_137(source_io_mem_137),
    .io_mem_138(source_io_mem_138),
    .io_mem_139(source_io_mem_139),
    .io_mem_140(source_io_mem_140),
    .io_mem_141(source_io_mem_141),
    .io_mem_142(source_io_mem_142),
    .io_mem_143(source_io_mem_143),
    .io_mem_144(source_io_mem_144),
    .io_mem_145(source_io_mem_145),
    .io_mem_146(source_io_mem_146),
    .io_mem_147(source_io_mem_147),
    .io_mem_148(source_io_mem_148),
    .io_mem_149(source_io_mem_149),
    .io_mem_150(source_io_mem_150),
    .io_mem_151(source_io_mem_151),
    .io_mem_152(source_io_mem_152),
    .io_mem_153(source_io_mem_153),
    .io_mem_154(source_io_mem_154),
    .io_mem_155(source_io_mem_155),
    .io_mem_156(source_io_mem_156),
    .io_mem_157(source_io_mem_157),
    .io_mem_158(source_io_mem_158),
    .io_mem_159(source_io_mem_159),
    .io_mem_160(source_io_mem_160),
    .io_mem_161(source_io_mem_161),
    .io_mem_162(source_io_mem_162),
    .io_mem_163(source_io_mem_163),
    .io_mem_164(source_io_mem_164),
    .io_mem_165(source_io_mem_165),
    .io_mem_166(source_io_mem_166),
    .io_mem_167(source_io_mem_167),
    .io_mem_168(source_io_mem_168),
    .io_mem_169(source_io_mem_169),
    .io_mem_170(source_io_mem_170),
    .io_mem_171(source_io_mem_171),
    .io_mem_172(source_io_mem_172),
    .io_mem_173(source_io_mem_173),
    .io_mem_174(source_io_mem_174),
    .io_mem_175(source_io_mem_175),
    .io_mem_176(source_io_mem_176),
    .io_mem_177(source_io_mem_177),
    .io_mem_178(source_io_mem_178),
    .io_mem_179(source_io_mem_179),
    .io_mem_180(source_io_mem_180),
    .io_mem_181(source_io_mem_181),
    .io_mem_182(source_io_mem_182),
    .io_mem_183(source_io_mem_183),
    .io_mem_184(source_io_mem_184),
    .io_mem_185(source_io_mem_185),
    .io_mem_186(source_io_mem_186),
    .io_mem_187(source_io_mem_187),
    .io_mem_188(source_io_mem_188),
    .io_mem_189(source_io_mem_189),
    .io_mem_190(source_io_mem_190),
    .io_mem_191(source_io_mem_191),
    .io_mem_192(source_io_mem_192),
    .io_mem_193(source_io_mem_193),
    .io_mem_194(source_io_mem_194),
    .io_mem_195(source_io_mem_195),
    .io_mem_196(source_io_mem_196),
    .io_mem_197(source_io_mem_197),
    .io_mem_198(source_io_mem_198),
    .io_mem_199(source_io_mem_199),
    .io_mem_200(source_io_mem_200),
    .io_mem_201(source_io_mem_201),
    .io_mem_202(source_io_mem_202),
    .io_mem_203(source_io_mem_203),
    .io_mem_204(source_io_mem_204),
    .io_mem_205(source_io_mem_205),
    .io_mem_206(source_io_mem_206),
    .io_mem_207(source_io_mem_207),
    .io_mem_208(source_io_mem_208),
    .io_mem_209(source_io_mem_209),
    .io_mem_210(source_io_mem_210),
    .io_mem_211(source_io_mem_211),
    .io_mem_212(source_io_mem_212),
    .io_mem_213(source_io_mem_213),
    .io_mem_214(source_io_mem_214),
    .io_mem_215(source_io_mem_215),
    .io_mem_216(source_io_mem_216),
    .io_mem_217(source_io_mem_217),
    .io_mem_218(source_io_mem_218),
    .io_mem_219(source_io_mem_219),
    .io_mem_220(source_io_mem_220),
    .io_mem_221(source_io_mem_221),
    .io_mem_222(source_io_mem_222),
    .io_mem_223(source_io_mem_223),
    .io_mem_224(source_io_mem_224),
    .io_mem_225(source_io_mem_225),
    .io_mem_226(source_io_mem_226),
    .io_mem_227(source_io_mem_227),
    .io_mem_228(source_io_mem_228),
    .io_mem_229(source_io_mem_229),
    .io_mem_230(source_io_mem_230),
    .io_mem_231(source_io_mem_231),
    .io_mem_232(source_io_mem_232),
    .io_mem_233(source_io_mem_233),
    .io_mem_234(source_io_mem_234),
    .io_mem_235(source_io_mem_235),
    .io_mem_236(source_io_mem_236),
    .io_mem_237(source_io_mem_237),
    .io_mem_238(source_io_mem_238),
    .io_mem_239(source_io_mem_239),
    .io_mem_240(source_io_mem_240),
    .io_mem_241(source_io_mem_241),
    .io_mem_242(source_io_mem_242),
    .io_mem_243(source_io_mem_243),
    .io_mem_244(source_io_mem_244),
    .io_mem_245(source_io_mem_245),
    .io_mem_246(source_io_mem_246),
    .io_mem_247(source_io_mem_247),
    .io_mem_248(source_io_mem_248),
    .io_mem_249(source_io_mem_249),
    .io_mem_250(source_io_mem_250),
    .io_mem_251(source_io_mem_251),
    .io_mem_252(source_io_mem_252),
    .io_mem_253(source_io_mem_253),
    .io_mem_254(source_io_mem_254),
    .io_mem_255(source_io_mem_255),
    .io_sink_reset_n(source_io_sink_reset_n),
    .io_ridx_valid(source_io_ridx_valid),
    .io_widx_valid(source_io_widx_valid)
  );
  AsyncQueueSink_1 sink ( // @[AsyncQueue.scala 156:22]
    .clock(sink_clock),
    .reset(sink_reset),
    .io_deq_ready(sink_io_deq_ready),
    .io_deq_valid(sink_io_deq_valid),
    .io_deq_bits(sink_io_deq_bits),
    .io_ridx(sink_io_ridx),
    .io_widx(sink_io_widx),
    .io_mem_0(sink_io_mem_0),
    .io_mem_1(sink_io_mem_1),
    .io_mem_2(sink_io_mem_2),
    .io_mem_3(sink_io_mem_3),
    .io_mem_4(sink_io_mem_4),
    .io_mem_5(sink_io_mem_5),
    .io_mem_6(sink_io_mem_6),
    .io_mem_7(sink_io_mem_7),
    .io_mem_8(sink_io_mem_8),
    .io_mem_9(sink_io_mem_9),
    .io_mem_10(sink_io_mem_10),
    .io_mem_11(sink_io_mem_11),
    .io_mem_12(sink_io_mem_12),
    .io_mem_13(sink_io_mem_13),
    .io_mem_14(sink_io_mem_14),
    .io_mem_15(sink_io_mem_15),
    .io_mem_16(sink_io_mem_16),
    .io_mem_17(sink_io_mem_17),
    .io_mem_18(sink_io_mem_18),
    .io_mem_19(sink_io_mem_19),
    .io_mem_20(sink_io_mem_20),
    .io_mem_21(sink_io_mem_21),
    .io_mem_22(sink_io_mem_22),
    .io_mem_23(sink_io_mem_23),
    .io_mem_24(sink_io_mem_24),
    .io_mem_25(sink_io_mem_25),
    .io_mem_26(sink_io_mem_26),
    .io_mem_27(sink_io_mem_27),
    .io_mem_28(sink_io_mem_28),
    .io_mem_29(sink_io_mem_29),
    .io_mem_30(sink_io_mem_30),
    .io_mem_31(sink_io_mem_31),
    .io_mem_32(sink_io_mem_32),
    .io_mem_33(sink_io_mem_33),
    .io_mem_34(sink_io_mem_34),
    .io_mem_35(sink_io_mem_35),
    .io_mem_36(sink_io_mem_36),
    .io_mem_37(sink_io_mem_37),
    .io_mem_38(sink_io_mem_38),
    .io_mem_39(sink_io_mem_39),
    .io_mem_40(sink_io_mem_40),
    .io_mem_41(sink_io_mem_41),
    .io_mem_42(sink_io_mem_42),
    .io_mem_43(sink_io_mem_43),
    .io_mem_44(sink_io_mem_44),
    .io_mem_45(sink_io_mem_45),
    .io_mem_46(sink_io_mem_46),
    .io_mem_47(sink_io_mem_47),
    .io_mem_48(sink_io_mem_48),
    .io_mem_49(sink_io_mem_49),
    .io_mem_50(sink_io_mem_50),
    .io_mem_51(sink_io_mem_51),
    .io_mem_52(sink_io_mem_52),
    .io_mem_53(sink_io_mem_53),
    .io_mem_54(sink_io_mem_54),
    .io_mem_55(sink_io_mem_55),
    .io_mem_56(sink_io_mem_56),
    .io_mem_57(sink_io_mem_57),
    .io_mem_58(sink_io_mem_58),
    .io_mem_59(sink_io_mem_59),
    .io_mem_60(sink_io_mem_60),
    .io_mem_61(sink_io_mem_61),
    .io_mem_62(sink_io_mem_62),
    .io_mem_63(sink_io_mem_63),
    .io_mem_64(sink_io_mem_64),
    .io_mem_65(sink_io_mem_65),
    .io_mem_66(sink_io_mem_66),
    .io_mem_67(sink_io_mem_67),
    .io_mem_68(sink_io_mem_68),
    .io_mem_69(sink_io_mem_69),
    .io_mem_70(sink_io_mem_70),
    .io_mem_71(sink_io_mem_71),
    .io_mem_72(sink_io_mem_72),
    .io_mem_73(sink_io_mem_73),
    .io_mem_74(sink_io_mem_74),
    .io_mem_75(sink_io_mem_75),
    .io_mem_76(sink_io_mem_76),
    .io_mem_77(sink_io_mem_77),
    .io_mem_78(sink_io_mem_78),
    .io_mem_79(sink_io_mem_79),
    .io_mem_80(sink_io_mem_80),
    .io_mem_81(sink_io_mem_81),
    .io_mem_82(sink_io_mem_82),
    .io_mem_83(sink_io_mem_83),
    .io_mem_84(sink_io_mem_84),
    .io_mem_85(sink_io_mem_85),
    .io_mem_86(sink_io_mem_86),
    .io_mem_87(sink_io_mem_87),
    .io_mem_88(sink_io_mem_88),
    .io_mem_89(sink_io_mem_89),
    .io_mem_90(sink_io_mem_90),
    .io_mem_91(sink_io_mem_91),
    .io_mem_92(sink_io_mem_92),
    .io_mem_93(sink_io_mem_93),
    .io_mem_94(sink_io_mem_94),
    .io_mem_95(sink_io_mem_95),
    .io_mem_96(sink_io_mem_96),
    .io_mem_97(sink_io_mem_97),
    .io_mem_98(sink_io_mem_98),
    .io_mem_99(sink_io_mem_99),
    .io_mem_100(sink_io_mem_100),
    .io_mem_101(sink_io_mem_101),
    .io_mem_102(sink_io_mem_102),
    .io_mem_103(sink_io_mem_103),
    .io_mem_104(sink_io_mem_104),
    .io_mem_105(sink_io_mem_105),
    .io_mem_106(sink_io_mem_106),
    .io_mem_107(sink_io_mem_107),
    .io_mem_108(sink_io_mem_108),
    .io_mem_109(sink_io_mem_109),
    .io_mem_110(sink_io_mem_110),
    .io_mem_111(sink_io_mem_111),
    .io_mem_112(sink_io_mem_112),
    .io_mem_113(sink_io_mem_113),
    .io_mem_114(sink_io_mem_114),
    .io_mem_115(sink_io_mem_115),
    .io_mem_116(sink_io_mem_116),
    .io_mem_117(sink_io_mem_117),
    .io_mem_118(sink_io_mem_118),
    .io_mem_119(sink_io_mem_119),
    .io_mem_120(sink_io_mem_120),
    .io_mem_121(sink_io_mem_121),
    .io_mem_122(sink_io_mem_122),
    .io_mem_123(sink_io_mem_123),
    .io_mem_124(sink_io_mem_124),
    .io_mem_125(sink_io_mem_125),
    .io_mem_126(sink_io_mem_126),
    .io_mem_127(sink_io_mem_127),
    .io_mem_128(sink_io_mem_128),
    .io_mem_129(sink_io_mem_129),
    .io_mem_130(sink_io_mem_130),
    .io_mem_131(sink_io_mem_131),
    .io_mem_132(sink_io_mem_132),
    .io_mem_133(sink_io_mem_133),
    .io_mem_134(sink_io_mem_134),
    .io_mem_135(sink_io_mem_135),
    .io_mem_136(sink_io_mem_136),
    .io_mem_137(sink_io_mem_137),
    .io_mem_138(sink_io_mem_138),
    .io_mem_139(sink_io_mem_139),
    .io_mem_140(sink_io_mem_140),
    .io_mem_141(sink_io_mem_141),
    .io_mem_142(sink_io_mem_142),
    .io_mem_143(sink_io_mem_143),
    .io_mem_144(sink_io_mem_144),
    .io_mem_145(sink_io_mem_145),
    .io_mem_146(sink_io_mem_146),
    .io_mem_147(sink_io_mem_147),
    .io_mem_148(sink_io_mem_148),
    .io_mem_149(sink_io_mem_149),
    .io_mem_150(sink_io_mem_150),
    .io_mem_151(sink_io_mem_151),
    .io_mem_152(sink_io_mem_152),
    .io_mem_153(sink_io_mem_153),
    .io_mem_154(sink_io_mem_154),
    .io_mem_155(sink_io_mem_155),
    .io_mem_156(sink_io_mem_156),
    .io_mem_157(sink_io_mem_157),
    .io_mem_158(sink_io_mem_158),
    .io_mem_159(sink_io_mem_159),
    .io_mem_160(sink_io_mem_160),
    .io_mem_161(sink_io_mem_161),
    .io_mem_162(sink_io_mem_162),
    .io_mem_163(sink_io_mem_163),
    .io_mem_164(sink_io_mem_164),
    .io_mem_165(sink_io_mem_165),
    .io_mem_166(sink_io_mem_166),
    .io_mem_167(sink_io_mem_167),
    .io_mem_168(sink_io_mem_168),
    .io_mem_169(sink_io_mem_169),
    .io_mem_170(sink_io_mem_170),
    .io_mem_171(sink_io_mem_171),
    .io_mem_172(sink_io_mem_172),
    .io_mem_173(sink_io_mem_173),
    .io_mem_174(sink_io_mem_174),
    .io_mem_175(sink_io_mem_175),
    .io_mem_176(sink_io_mem_176),
    .io_mem_177(sink_io_mem_177),
    .io_mem_178(sink_io_mem_178),
    .io_mem_179(sink_io_mem_179),
    .io_mem_180(sink_io_mem_180),
    .io_mem_181(sink_io_mem_181),
    .io_mem_182(sink_io_mem_182),
    .io_mem_183(sink_io_mem_183),
    .io_mem_184(sink_io_mem_184),
    .io_mem_185(sink_io_mem_185),
    .io_mem_186(sink_io_mem_186),
    .io_mem_187(sink_io_mem_187),
    .io_mem_188(sink_io_mem_188),
    .io_mem_189(sink_io_mem_189),
    .io_mem_190(sink_io_mem_190),
    .io_mem_191(sink_io_mem_191),
    .io_mem_192(sink_io_mem_192),
    .io_mem_193(sink_io_mem_193),
    .io_mem_194(sink_io_mem_194),
    .io_mem_195(sink_io_mem_195),
    .io_mem_196(sink_io_mem_196),
    .io_mem_197(sink_io_mem_197),
    .io_mem_198(sink_io_mem_198),
    .io_mem_199(sink_io_mem_199),
    .io_mem_200(sink_io_mem_200),
    .io_mem_201(sink_io_mem_201),
    .io_mem_202(sink_io_mem_202),
    .io_mem_203(sink_io_mem_203),
    .io_mem_204(sink_io_mem_204),
    .io_mem_205(sink_io_mem_205),
    .io_mem_206(sink_io_mem_206),
    .io_mem_207(sink_io_mem_207),
    .io_mem_208(sink_io_mem_208),
    .io_mem_209(sink_io_mem_209),
    .io_mem_210(sink_io_mem_210),
    .io_mem_211(sink_io_mem_211),
    .io_mem_212(sink_io_mem_212),
    .io_mem_213(sink_io_mem_213),
    .io_mem_214(sink_io_mem_214),
    .io_mem_215(sink_io_mem_215),
    .io_mem_216(sink_io_mem_216),
    .io_mem_217(sink_io_mem_217),
    .io_mem_218(sink_io_mem_218),
    .io_mem_219(sink_io_mem_219),
    .io_mem_220(sink_io_mem_220),
    .io_mem_221(sink_io_mem_221),
    .io_mem_222(sink_io_mem_222),
    .io_mem_223(sink_io_mem_223),
    .io_mem_224(sink_io_mem_224),
    .io_mem_225(sink_io_mem_225),
    .io_mem_226(sink_io_mem_226),
    .io_mem_227(sink_io_mem_227),
    .io_mem_228(sink_io_mem_228),
    .io_mem_229(sink_io_mem_229),
    .io_mem_230(sink_io_mem_230),
    .io_mem_231(sink_io_mem_231),
    .io_mem_232(sink_io_mem_232),
    .io_mem_233(sink_io_mem_233),
    .io_mem_234(sink_io_mem_234),
    .io_mem_235(sink_io_mem_235),
    .io_mem_236(sink_io_mem_236),
    .io_mem_237(sink_io_mem_237),
    .io_mem_238(sink_io_mem_238),
    .io_mem_239(sink_io_mem_239),
    .io_mem_240(sink_io_mem_240),
    .io_mem_241(sink_io_mem_241),
    .io_mem_242(sink_io_mem_242),
    .io_mem_243(sink_io_mem_243),
    .io_mem_244(sink_io_mem_244),
    .io_mem_245(sink_io_mem_245),
    .io_mem_246(sink_io_mem_246),
    .io_mem_247(sink_io_mem_247),
    .io_mem_248(sink_io_mem_248),
    .io_mem_249(sink_io_mem_249),
    .io_mem_250(sink_io_mem_250),
    .io_mem_251(sink_io_mem_251),
    .io_mem_252(sink_io_mem_252),
    .io_mem_253(sink_io_mem_253),
    .io_mem_254(sink_io_mem_254),
    .io_mem_255(sink_io_mem_255),
    .io_source_reset_n(sink_io_source_reset_n),
    .io_ridx_valid(sink_io_ridx_valid),
    .io_widx_valid(sink_io_widx_valid)
  );
  assign io_enq_ready = source_io_enq_ready;
  assign io_deq_valid = sink_io_deq_valid;
  assign io_deq_bits = sink_io_deq_bits;
  assign source_clock = io_enq_clock;
  assign source_reset = 1'h0;
  assign source_io_enq_valid = io_enq_valid;
  assign source_io_enq_bits = io_enq_bits;
  assign source_io_ridx = sink_io_ridx;
  assign source_io_sink_reset_n = 1'h1;
  assign source_io_ridx_valid = sink_io_ridx_valid;
  assign sink_clock = io_deq_clock;
  assign sink_reset = 1'h0;
  assign sink_io_deq_ready = io_deq_ready;
  assign sink_io_widx = source_io_widx;
  assign sink_io_mem_0 = source_io_mem_0;
  assign sink_io_mem_1 = source_io_mem_1;
  assign sink_io_mem_2 = source_io_mem_2;
  assign sink_io_mem_3 = source_io_mem_3;
  assign sink_io_mem_4 = source_io_mem_4;
  assign sink_io_mem_5 = source_io_mem_5;
  assign sink_io_mem_6 = source_io_mem_6;
  assign sink_io_mem_7 = source_io_mem_7;
  assign sink_io_mem_8 = source_io_mem_8;
  assign sink_io_mem_9 = source_io_mem_9;
  assign sink_io_mem_10 = source_io_mem_10;
  assign sink_io_mem_11 = source_io_mem_11;
  assign sink_io_mem_12 = source_io_mem_12;
  assign sink_io_mem_13 = source_io_mem_13;
  assign sink_io_mem_14 = source_io_mem_14;
  assign sink_io_mem_15 = source_io_mem_15;
  assign sink_io_mem_16 = source_io_mem_16;
  assign sink_io_mem_17 = source_io_mem_17;
  assign sink_io_mem_18 = source_io_mem_18;
  assign sink_io_mem_19 = source_io_mem_19;
  assign sink_io_mem_20 = source_io_mem_20;
  assign sink_io_mem_21 = source_io_mem_21;
  assign sink_io_mem_22 = source_io_mem_22;
  assign sink_io_mem_23 = source_io_mem_23;
  assign sink_io_mem_24 = source_io_mem_24;
  assign sink_io_mem_25 = source_io_mem_25;
  assign sink_io_mem_26 = source_io_mem_26;
  assign sink_io_mem_27 = source_io_mem_27;
  assign sink_io_mem_28 = source_io_mem_28;
  assign sink_io_mem_29 = source_io_mem_29;
  assign sink_io_mem_30 = source_io_mem_30;
  assign sink_io_mem_31 = source_io_mem_31;
  assign sink_io_mem_32 = source_io_mem_32;
  assign sink_io_mem_33 = source_io_mem_33;
  assign sink_io_mem_34 = source_io_mem_34;
  assign sink_io_mem_35 = source_io_mem_35;
  assign sink_io_mem_36 = source_io_mem_36;
  assign sink_io_mem_37 = source_io_mem_37;
  assign sink_io_mem_38 = source_io_mem_38;
  assign sink_io_mem_39 = source_io_mem_39;
  assign sink_io_mem_40 = source_io_mem_40;
  assign sink_io_mem_41 = source_io_mem_41;
  assign sink_io_mem_42 = source_io_mem_42;
  assign sink_io_mem_43 = source_io_mem_43;
  assign sink_io_mem_44 = source_io_mem_44;
  assign sink_io_mem_45 = source_io_mem_45;
  assign sink_io_mem_46 = source_io_mem_46;
  assign sink_io_mem_47 = source_io_mem_47;
  assign sink_io_mem_48 = source_io_mem_48;
  assign sink_io_mem_49 = source_io_mem_49;
  assign sink_io_mem_50 = source_io_mem_50;
  assign sink_io_mem_51 = source_io_mem_51;
  assign sink_io_mem_52 = source_io_mem_52;
  assign sink_io_mem_53 = source_io_mem_53;
  assign sink_io_mem_54 = source_io_mem_54;
  assign sink_io_mem_55 = source_io_mem_55;
  assign sink_io_mem_56 = source_io_mem_56;
  assign sink_io_mem_57 = source_io_mem_57;
  assign sink_io_mem_58 = source_io_mem_58;
  assign sink_io_mem_59 = source_io_mem_59;
  assign sink_io_mem_60 = source_io_mem_60;
  assign sink_io_mem_61 = source_io_mem_61;
  assign sink_io_mem_62 = source_io_mem_62;
  assign sink_io_mem_63 = source_io_mem_63;
  assign sink_io_mem_64 = source_io_mem_64;
  assign sink_io_mem_65 = source_io_mem_65;
  assign sink_io_mem_66 = source_io_mem_66;
  assign sink_io_mem_67 = source_io_mem_67;
  assign sink_io_mem_68 = source_io_mem_68;
  assign sink_io_mem_69 = source_io_mem_69;
  assign sink_io_mem_70 = source_io_mem_70;
  assign sink_io_mem_71 = source_io_mem_71;
  assign sink_io_mem_72 = source_io_mem_72;
  assign sink_io_mem_73 = source_io_mem_73;
  assign sink_io_mem_74 = source_io_mem_74;
  assign sink_io_mem_75 = source_io_mem_75;
  assign sink_io_mem_76 = source_io_mem_76;
  assign sink_io_mem_77 = source_io_mem_77;
  assign sink_io_mem_78 = source_io_mem_78;
  assign sink_io_mem_79 = source_io_mem_79;
  assign sink_io_mem_80 = source_io_mem_80;
  assign sink_io_mem_81 = source_io_mem_81;
  assign sink_io_mem_82 = source_io_mem_82;
  assign sink_io_mem_83 = source_io_mem_83;
  assign sink_io_mem_84 = source_io_mem_84;
  assign sink_io_mem_85 = source_io_mem_85;
  assign sink_io_mem_86 = source_io_mem_86;
  assign sink_io_mem_87 = source_io_mem_87;
  assign sink_io_mem_88 = source_io_mem_88;
  assign sink_io_mem_89 = source_io_mem_89;
  assign sink_io_mem_90 = source_io_mem_90;
  assign sink_io_mem_91 = source_io_mem_91;
  assign sink_io_mem_92 = source_io_mem_92;
  assign sink_io_mem_93 = source_io_mem_93;
  assign sink_io_mem_94 = source_io_mem_94;
  assign sink_io_mem_95 = source_io_mem_95;
  assign sink_io_mem_96 = source_io_mem_96;
  assign sink_io_mem_97 = source_io_mem_97;
  assign sink_io_mem_98 = source_io_mem_98;
  assign sink_io_mem_99 = source_io_mem_99;
  assign sink_io_mem_100 = source_io_mem_100;
  assign sink_io_mem_101 = source_io_mem_101;
  assign sink_io_mem_102 = source_io_mem_102;
  assign sink_io_mem_103 = source_io_mem_103;
  assign sink_io_mem_104 = source_io_mem_104;
  assign sink_io_mem_105 = source_io_mem_105;
  assign sink_io_mem_106 = source_io_mem_106;
  assign sink_io_mem_107 = source_io_mem_107;
  assign sink_io_mem_108 = source_io_mem_108;
  assign sink_io_mem_109 = source_io_mem_109;
  assign sink_io_mem_110 = source_io_mem_110;
  assign sink_io_mem_111 = source_io_mem_111;
  assign sink_io_mem_112 = source_io_mem_112;
  assign sink_io_mem_113 = source_io_mem_113;
  assign sink_io_mem_114 = source_io_mem_114;
  assign sink_io_mem_115 = source_io_mem_115;
  assign sink_io_mem_116 = source_io_mem_116;
  assign sink_io_mem_117 = source_io_mem_117;
  assign sink_io_mem_118 = source_io_mem_118;
  assign sink_io_mem_119 = source_io_mem_119;
  assign sink_io_mem_120 = source_io_mem_120;
  assign sink_io_mem_121 = source_io_mem_121;
  assign sink_io_mem_122 = source_io_mem_122;
  assign sink_io_mem_123 = source_io_mem_123;
  assign sink_io_mem_124 = source_io_mem_124;
  assign sink_io_mem_125 = source_io_mem_125;
  assign sink_io_mem_126 = source_io_mem_126;
  assign sink_io_mem_127 = source_io_mem_127;
  assign sink_io_mem_128 = source_io_mem_128;
  assign sink_io_mem_129 = source_io_mem_129;
  assign sink_io_mem_130 = source_io_mem_130;
  assign sink_io_mem_131 = source_io_mem_131;
  assign sink_io_mem_132 = source_io_mem_132;
  assign sink_io_mem_133 = source_io_mem_133;
  assign sink_io_mem_134 = source_io_mem_134;
  assign sink_io_mem_135 = source_io_mem_135;
  assign sink_io_mem_136 = source_io_mem_136;
  assign sink_io_mem_137 = source_io_mem_137;
  assign sink_io_mem_138 = source_io_mem_138;
  assign sink_io_mem_139 = source_io_mem_139;
  assign sink_io_mem_140 = source_io_mem_140;
  assign sink_io_mem_141 = source_io_mem_141;
  assign sink_io_mem_142 = source_io_mem_142;
  assign sink_io_mem_143 = source_io_mem_143;
  assign sink_io_mem_144 = source_io_mem_144;
  assign sink_io_mem_145 = source_io_mem_145;
  assign sink_io_mem_146 = source_io_mem_146;
  assign sink_io_mem_147 = source_io_mem_147;
  assign sink_io_mem_148 = source_io_mem_148;
  assign sink_io_mem_149 = source_io_mem_149;
  assign sink_io_mem_150 = source_io_mem_150;
  assign sink_io_mem_151 = source_io_mem_151;
  assign sink_io_mem_152 = source_io_mem_152;
  assign sink_io_mem_153 = source_io_mem_153;
  assign sink_io_mem_154 = source_io_mem_154;
  assign sink_io_mem_155 = source_io_mem_155;
  assign sink_io_mem_156 = source_io_mem_156;
  assign sink_io_mem_157 = source_io_mem_157;
  assign sink_io_mem_158 = source_io_mem_158;
  assign sink_io_mem_159 = source_io_mem_159;
  assign sink_io_mem_160 = source_io_mem_160;
  assign sink_io_mem_161 = source_io_mem_161;
  assign sink_io_mem_162 = source_io_mem_162;
  assign sink_io_mem_163 = source_io_mem_163;
  assign sink_io_mem_164 = source_io_mem_164;
  assign sink_io_mem_165 = source_io_mem_165;
  assign sink_io_mem_166 = source_io_mem_166;
  assign sink_io_mem_167 = source_io_mem_167;
  assign sink_io_mem_168 = source_io_mem_168;
  assign sink_io_mem_169 = source_io_mem_169;
  assign sink_io_mem_170 = source_io_mem_170;
  assign sink_io_mem_171 = source_io_mem_171;
  assign sink_io_mem_172 = source_io_mem_172;
  assign sink_io_mem_173 = source_io_mem_173;
  assign sink_io_mem_174 = source_io_mem_174;
  assign sink_io_mem_175 = source_io_mem_175;
  assign sink_io_mem_176 = source_io_mem_176;
  assign sink_io_mem_177 = source_io_mem_177;
  assign sink_io_mem_178 = source_io_mem_178;
  assign sink_io_mem_179 = source_io_mem_179;
  assign sink_io_mem_180 = source_io_mem_180;
  assign sink_io_mem_181 = source_io_mem_181;
  assign sink_io_mem_182 = source_io_mem_182;
  assign sink_io_mem_183 = source_io_mem_183;
  assign sink_io_mem_184 = source_io_mem_184;
  assign sink_io_mem_185 = source_io_mem_185;
  assign sink_io_mem_186 = source_io_mem_186;
  assign sink_io_mem_187 = source_io_mem_187;
  assign sink_io_mem_188 = source_io_mem_188;
  assign sink_io_mem_189 = source_io_mem_189;
  assign sink_io_mem_190 = source_io_mem_190;
  assign sink_io_mem_191 = source_io_mem_191;
  assign sink_io_mem_192 = source_io_mem_192;
  assign sink_io_mem_193 = source_io_mem_193;
  assign sink_io_mem_194 = source_io_mem_194;
  assign sink_io_mem_195 = source_io_mem_195;
  assign sink_io_mem_196 = source_io_mem_196;
  assign sink_io_mem_197 = source_io_mem_197;
  assign sink_io_mem_198 = source_io_mem_198;
  assign sink_io_mem_199 = source_io_mem_199;
  assign sink_io_mem_200 = source_io_mem_200;
  assign sink_io_mem_201 = source_io_mem_201;
  assign sink_io_mem_202 = source_io_mem_202;
  assign sink_io_mem_203 = source_io_mem_203;
  assign sink_io_mem_204 = source_io_mem_204;
  assign sink_io_mem_205 = source_io_mem_205;
  assign sink_io_mem_206 = source_io_mem_206;
  assign sink_io_mem_207 = source_io_mem_207;
  assign sink_io_mem_208 = source_io_mem_208;
  assign sink_io_mem_209 = source_io_mem_209;
  assign sink_io_mem_210 = source_io_mem_210;
  assign sink_io_mem_211 = source_io_mem_211;
  assign sink_io_mem_212 = source_io_mem_212;
  assign sink_io_mem_213 = source_io_mem_213;
  assign sink_io_mem_214 = source_io_mem_214;
  assign sink_io_mem_215 = source_io_mem_215;
  assign sink_io_mem_216 = source_io_mem_216;
  assign sink_io_mem_217 = source_io_mem_217;
  assign sink_io_mem_218 = source_io_mem_218;
  assign sink_io_mem_219 = source_io_mem_219;
  assign sink_io_mem_220 = source_io_mem_220;
  assign sink_io_mem_221 = source_io_mem_221;
  assign sink_io_mem_222 = source_io_mem_222;
  assign sink_io_mem_223 = source_io_mem_223;
  assign sink_io_mem_224 = source_io_mem_224;
  assign sink_io_mem_225 = source_io_mem_225;
  assign sink_io_mem_226 = source_io_mem_226;
  assign sink_io_mem_227 = source_io_mem_227;
  assign sink_io_mem_228 = source_io_mem_228;
  assign sink_io_mem_229 = source_io_mem_229;
  assign sink_io_mem_230 = source_io_mem_230;
  assign sink_io_mem_231 = source_io_mem_231;
  assign sink_io_mem_232 = source_io_mem_232;
  assign sink_io_mem_233 = source_io_mem_233;
  assign sink_io_mem_234 = source_io_mem_234;
  assign sink_io_mem_235 = source_io_mem_235;
  assign sink_io_mem_236 = source_io_mem_236;
  assign sink_io_mem_237 = source_io_mem_237;
  assign sink_io_mem_238 = source_io_mem_238;
  assign sink_io_mem_239 = source_io_mem_239;
  assign sink_io_mem_240 = source_io_mem_240;
  assign sink_io_mem_241 = source_io_mem_241;
  assign sink_io_mem_242 = source_io_mem_242;
  assign sink_io_mem_243 = source_io_mem_243;
  assign sink_io_mem_244 = source_io_mem_244;
  assign sink_io_mem_245 = source_io_mem_245;
  assign sink_io_mem_246 = source_io_mem_246;
  assign sink_io_mem_247 = source_io_mem_247;
  assign sink_io_mem_248 = source_io_mem_248;
  assign sink_io_mem_249 = source_io_mem_249;
  assign sink_io_mem_250 = source_io_mem_250;
  assign sink_io_mem_251 = source_io_mem_251;
  assign sink_io_mem_252 = source_io_mem_252;
  assign sink_io_mem_253 = source_io_mem_253;
  assign sink_io_mem_254 = source_io_mem_254;
  assign sink_io_mem_255 = source_io_mem_255;
  assign sink_io_source_reset_n = 1'h1;
  assign sink_io_widx_valid = source_io_widx_valid;
endmodule
module PDATop(
  input         io_ARM_Switch_i,
  input  [31:0] io_ARM_AA_i,
  input  [23:0] io_ARM_CRC_Seed_i,
  input  [6:0]  io_ARM_DeWhite_Seed_i,
  input         io_ARM_Data_o_ready,
  output        io_ARM_Data_o_valid,
  output [7:0]  io_ARM_Data_o_bits,
  input         io_ARM_Length_o_ready,
  output        io_ARM_Length_o_valid,
  output [7:0]  io_ARM_Length_o_bits,
  input         io_ARM_Flag_AA_o_ready,
  output        io_ARM_Flag_AA_o_valid,
  output        io_ARM_Flag_AA_o_bits,
  input         io_ARM_Flag_CRC_o_ready,
  output        io_ARM_Flag_CRC_o_valid,
  output        io_ARM_Flag_CRC_o_bits,
  input         io_CDR_recovered_clk,
  input         io_CDR_recovered_data,
  output        io_ARM_data_i_ready,
  input         io_ARM_data_i_valid,
  input         io_ARM_data_i_bits,
  input         io_choose_data_src,
  input         io_clk_CDR,
  input         io_reset_CDR,
  input         io_clk_PDA,
  input         io_clk_ARM
);
  wire  ble_packetdisassembler_clock; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_reset; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_DMA_Switch_i; // @[PDATop.scala 69:21]
  wire [31:0] ble_packetdisassembler_io_REG_AA_i; // @[PDATop.scala 69:21]
  wire [23:0] ble_packetdisassembler_io_REG_CRC_Seed_i; // @[PDATop.scala 69:21]
  wire [6:0] ble_packetdisassembler_io_REG_DeWhite_Seed_i; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_DMA_Data_o_ready; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_DMA_Data_o_valid; // @[PDATop.scala 69:21]
  wire [7:0] ble_packetdisassembler_io_DMA_Data_o_bits; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_DMA_Length_o_ready; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_DMA_Length_o_valid; // @[PDATop.scala 69:21]
  wire [7:0] ble_packetdisassembler_io_DMA_Length_o_bits; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_DMA_Flag_AA_o_ready; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_DMA_Flag_AA_o_valid; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_DMA_Flag_AA_o_bits; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_DMA_Flag_CRC_o_ready; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_DMA_Flag_CRC_o_valid; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_DMA_Flag_CRC_o_bits; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_AFIFO_Data_i_ready; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_AFIFO_Data_i_valid; // @[PDATop.scala 69:21]
  wire  ble_packetdisassembler_io_AFIFO_Data_i_bits; // @[PDATop.scala 69:21]
  wire  AsyncQueue_io_enq_clock; // @[PDATop.scala 80:27]
  wire  AsyncQueue_io_enq_ready; // @[PDATop.scala 80:27]
  wire  AsyncQueue_io_enq_valid; // @[PDATop.scala 80:27]
  wire  AsyncQueue_io_enq_bits; // @[PDATop.scala 80:27]
  wire  AsyncQueue_io_deq_clock; // @[PDATop.scala 80:27]
  wire  AsyncQueue_io_deq_ready; // @[PDATop.scala 80:27]
  wire  AsyncQueue_io_deq_valid; // @[PDATop.scala 80:27]
  wire  AsyncQueue_io_deq_bits; // @[PDATop.scala 80:27]
  wire  AsyncQueue_1_io_enq_clock; // @[PDATop.scala 101:26]
  wire  AsyncQueue_1_io_enq_ready; // @[PDATop.scala 101:26]
  wire  AsyncQueue_1_io_enq_valid; // @[PDATop.scala 101:26]
  wire [7:0] AsyncQueue_1_io_enq_bits; // @[PDATop.scala 101:26]
  wire  AsyncQueue_1_io_deq_clock; // @[PDATop.scala 101:26]
  wire  AsyncQueue_1_io_deq_ready; // @[PDATop.scala 101:26]
  wire  AsyncQueue_1_io_deq_valid; // @[PDATop.scala 101:26]
  wire [7:0] AsyncQueue_1_io_deq_bits; // @[PDATop.scala 101:26]
  wire  AsyncQueue_2_io_enq_clock; // @[PDATop.scala 101:26]
  wire  AsyncQueue_2_io_enq_ready; // @[PDATop.scala 101:26]
  wire  AsyncQueue_2_io_enq_valid; // @[PDATop.scala 101:26]
  wire [7:0] AsyncQueue_2_io_enq_bits; // @[PDATop.scala 101:26]
  wire  AsyncQueue_2_io_deq_clock; // @[PDATop.scala 101:26]
  wire  AsyncQueue_2_io_deq_ready; // @[PDATop.scala 101:26]
  wire  AsyncQueue_2_io_deq_valid; // @[PDATop.scala 101:26]
  wire [7:0] AsyncQueue_2_io_deq_bits; // @[PDATop.scala 101:26]
  wire  AsyncQueue_3_io_enq_clock; // @[PDATop.scala 101:26]
  wire  AsyncQueue_3_io_enq_ready; // @[PDATop.scala 101:26]
  wire  AsyncQueue_3_io_enq_valid; // @[PDATop.scala 101:26]
  wire  AsyncQueue_3_io_enq_bits; // @[PDATop.scala 101:26]
  wire  AsyncQueue_3_io_deq_clock; // @[PDATop.scala 101:26]
  wire  AsyncQueue_3_io_deq_ready; // @[PDATop.scala 101:26]
  wire  AsyncQueue_3_io_deq_valid; // @[PDATop.scala 101:26]
  wire  AsyncQueue_3_io_deq_bits; // @[PDATop.scala 101:26]
  wire  AsyncQueue_4_io_enq_clock; // @[PDATop.scala 101:26]
  wire  AsyncQueue_4_io_enq_ready; // @[PDATop.scala 101:26]
  wire  AsyncQueue_4_io_enq_valid; // @[PDATop.scala 101:26]
  wire  AsyncQueue_4_io_enq_bits; // @[PDATop.scala 101:26]
  wire  AsyncQueue_4_io_deq_clock; // @[PDATop.scala 101:26]
  wire  AsyncQueue_4_io_deq_ready; // @[PDATop.scala 101:26]
  wire  AsyncQueue_4_io_deq_valid; // @[PDATop.scala 101:26]
  wire  AsyncQueue_4_io_deq_bits; // @[PDATop.scala 101:26]
  wire  _T_40_bits; // @[PDATop.scala 77:28]
  wire  _T_48; // @[PDATop.scala 94:36]
  wire  _T_40_valid; // @[PDATop.scala 77:28]
  wire  _T_49; // @[PDATop.scala 95:37]
  wire  _T_40_ready; // @[PDATop.scala 77:28]
  ble_packetdisassembler ble_packetdisassembler ( // @[PDATop.scala 69:21]
    .clock(ble_packetdisassembler_clock),
    .reset(ble_packetdisassembler_reset),
    .io_DMA_Switch_i(ble_packetdisassembler_io_DMA_Switch_i),
    .io_REG_AA_i(ble_packetdisassembler_io_REG_AA_i),
    .io_REG_CRC_Seed_i(ble_packetdisassembler_io_REG_CRC_Seed_i),
    .io_REG_DeWhite_Seed_i(ble_packetdisassembler_io_REG_DeWhite_Seed_i),
    .io_DMA_Data_o_ready(ble_packetdisassembler_io_DMA_Data_o_ready),
    .io_DMA_Data_o_valid(ble_packetdisassembler_io_DMA_Data_o_valid),
    .io_DMA_Data_o_bits(ble_packetdisassembler_io_DMA_Data_o_bits),
    .io_DMA_Length_o_ready(ble_packetdisassembler_io_DMA_Length_o_ready),
    .io_DMA_Length_o_valid(ble_packetdisassembler_io_DMA_Length_o_valid),
    .io_DMA_Length_o_bits(ble_packetdisassembler_io_DMA_Length_o_bits),
    .io_DMA_Flag_AA_o_ready(ble_packetdisassembler_io_DMA_Flag_AA_o_ready),
    .io_DMA_Flag_AA_o_valid(ble_packetdisassembler_io_DMA_Flag_AA_o_valid),
    .io_DMA_Flag_AA_o_bits(ble_packetdisassembler_io_DMA_Flag_AA_o_bits),
    .io_DMA_Flag_CRC_o_ready(ble_packetdisassembler_io_DMA_Flag_CRC_o_ready),
    .io_DMA_Flag_CRC_o_valid(ble_packetdisassembler_io_DMA_Flag_CRC_o_valid),
    .io_DMA_Flag_CRC_o_bits(ble_packetdisassembler_io_DMA_Flag_CRC_o_bits),
    .io_AFIFO_Data_i_ready(ble_packetdisassembler_io_AFIFO_Data_i_ready),
    .io_AFIFO_Data_i_valid(ble_packetdisassembler_io_AFIFO_Data_i_valid),
    .io_AFIFO_Data_i_bits(ble_packetdisassembler_io_AFIFO_Data_i_bits)
  );
  AsyncQueue AsyncQueue ( // @[PDATop.scala 80:27]
    .io_enq_clock(AsyncQueue_io_enq_clock),
    .io_enq_ready(AsyncQueue_io_enq_ready),
    .io_enq_valid(AsyncQueue_io_enq_valid),
    .io_enq_bits(AsyncQueue_io_enq_bits),
    .io_deq_clock(AsyncQueue_io_deq_clock),
    .io_deq_ready(AsyncQueue_io_deq_ready),
    .io_deq_valid(AsyncQueue_io_deq_valid),
    .io_deq_bits(AsyncQueue_io_deq_bits)
  );
  AsyncQueue_1 AsyncQueue_1 ( // @[PDATop.scala 101:26]
    .io_enq_clock(AsyncQueue_1_io_enq_clock),
    .io_enq_ready(AsyncQueue_1_io_enq_ready),
    .io_enq_valid(AsyncQueue_1_io_enq_valid),
    .io_enq_bits(AsyncQueue_1_io_enq_bits),
    .io_deq_clock(AsyncQueue_1_io_deq_clock),
    .io_deq_ready(AsyncQueue_1_io_deq_ready),
    .io_deq_valid(AsyncQueue_1_io_deq_valid),
    .io_deq_bits(AsyncQueue_1_io_deq_bits)
  );
  AsyncQueue_1 AsyncQueue_2 ( // @[PDATop.scala 101:26]
    .io_enq_clock(AsyncQueue_2_io_enq_clock),
    .io_enq_ready(AsyncQueue_2_io_enq_ready),
    .io_enq_valid(AsyncQueue_2_io_enq_valid),
    .io_enq_bits(AsyncQueue_2_io_enq_bits),
    .io_deq_clock(AsyncQueue_2_io_deq_clock),
    .io_deq_ready(AsyncQueue_2_io_deq_ready),
    .io_deq_valid(AsyncQueue_2_io_deq_valid),
    .io_deq_bits(AsyncQueue_2_io_deq_bits)
  );
  AsyncQueue AsyncQueue_3 ( // @[PDATop.scala 101:26]
    .io_enq_clock(AsyncQueue_3_io_enq_clock),
    .io_enq_ready(AsyncQueue_3_io_enq_ready),
    .io_enq_valid(AsyncQueue_3_io_enq_valid),
    .io_enq_bits(AsyncQueue_3_io_enq_bits),
    .io_deq_clock(AsyncQueue_3_io_deq_clock),
    .io_deq_ready(AsyncQueue_3_io_deq_ready),
    .io_deq_valid(AsyncQueue_3_io_deq_valid),
    .io_deq_bits(AsyncQueue_3_io_deq_bits)
  );
  AsyncQueue AsyncQueue_4 ( // @[PDATop.scala 101:26]
    .io_enq_clock(AsyncQueue_4_io_enq_clock),
    .io_enq_ready(AsyncQueue_4_io_enq_ready),
    .io_enq_valid(AsyncQueue_4_io_enq_valid),
    .io_enq_bits(AsyncQueue_4_io_enq_bits),
    .io_deq_clock(AsyncQueue_4_io_deq_clock),
    .io_deq_ready(AsyncQueue_4_io_deq_ready),
    .io_deq_valid(AsyncQueue_4_io_deq_valid),
    .io_deq_bits(AsyncQueue_4_io_deq_bits)
  );
  assign _T_40_bits = AsyncQueue_io_deq_bits; // @[PDATop.scala 77:28]
  assign _T_48 = io_choose_data_src ? io_ARM_data_i_bits : _T_40_bits; // @[PDATop.scala 94:36]
  assign _T_40_valid = AsyncQueue_io_deq_valid; // @[PDATop.scala 77:28]
  assign _T_49 = io_choose_data_src ? io_ARM_data_i_valid : _T_40_valid; // @[PDATop.scala 95:37]
  assign _T_40_ready = ble_packetdisassembler_io_AFIFO_Data_i_ready; // @[PDATop.scala 77:28]
  assign io_ARM_Data_o_valid = AsyncQueue_1_io_deq_valid;
  assign io_ARM_Data_o_bits = AsyncQueue_1_io_deq_bits;
  assign io_ARM_Length_o_valid = AsyncQueue_2_io_deq_valid;
  assign io_ARM_Length_o_bits = AsyncQueue_2_io_deq_bits;
  assign io_ARM_Flag_AA_o_valid = AsyncQueue_3_io_deq_valid;
  assign io_ARM_Flag_AA_o_bits = AsyncQueue_3_io_deq_bits;
  assign io_ARM_Flag_CRC_o_valid = AsyncQueue_4_io_deq_valid;
  assign io_ARM_Flag_CRC_o_bits = AsyncQueue_4_io_deq_bits;
  assign io_ARM_data_i_ready = ble_packetdisassembler_io_AFIFO_Data_i_ready;
  assign ble_packetdisassembler_clock = io_clk_CDR;
  assign ble_packetdisassembler_reset = io_reset_CDR;
  assign ble_packetdisassembler_io_DMA_Switch_i = io_ARM_Switch_i;
  assign ble_packetdisassembler_io_REG_AA_i = io_ARM_AA_i;
  assign ble_packetdisassembler_io_REG_CRC_Seed_i = io_ARM_CRC_Seed_i;
  assign ble_packetdisassembler_io_REG_DeWhite_Seed_i = io_ARM_DeWhite_Seed_i;
  assign ble_packetdisassembler_io_DMA_Data_o_ready = AsyncQueue_1_io_enq_ready;
  assign ble_packetdisassembler_io_DMA_Length_o_ready = AsyncQueue_2_io_enq_ready;
  assign ble_packetdisassembler_io_DMA_Flag_AA_o_ready = AsyncQueue_3_io_enq_ready;
  assign ble_packetdisassembler_io_DMA_Flag_CRC_o_ready = AsyncQueue_4_io_enq_ready;
  assign ble_packetdisassembler_io_AFIFO_Data_i_valid = _T_49;
  assign ble_packetdisassembler_io_AFIFO_Data_i_bits = _T_48;
  assign AsyncQueue_io_enq_clock = io_clk_CDR;
  assign AsyncQueue_io_enq_valid = io_CDR_recovered_clk;
  assign AsyncQueue_io_enq_bits = io_CDR_recovered_data;
  assign AsyncQueue_io_deq_clock = io_clk_PDA;
  assign AsyncQueue_io_deq_ready = _T_40_ready;
  assign AsyncQueue_1_io_enq_clock = io_clk_PDA;
  assign AsyncQueue_1_io_enq_valid = ble_packetdisassembler_io_DMA_Data_o_valid;
  assign AsyncQueue_1_io_enq_bits = ble_packetdisassembler_io_DMA_Data_o_bits;
  assign AsyncQueue_1_io_deq_clock = io_clk_ARM;
  assign AsyncQueue_1_io_deq_ready = io_ARM_Data_o_ready;
  assign AsyncQueue_2_io_enq_clock = io_clk_PDA;
  assign AsyncQueue_2_io_enq_valid = ble_packetdisassembler_io_DMA_Length_o_valid;
  assign AsyncQueue_2_io_enq_bits = ble_packetdisassembler_io_DMA_Length_o_bits;
  assign AsyncQueue_2_io_deq_clock = io_clk_ARM;
  assign AsyncQueue_2_io_deq_ready = io_ARM_Length_o_ready;
  assign AsyncQueue_3_io_enq_clock = io_clk_PDA;
  assign AsyncQueue_3_io_enq_valid = ble_packetdisassembler_io_DMA_Flag_AA_o_valid;
  assign AsyncQueue_3_io_enq_bits = ble_packetdisassembler_io_DMA_Flag_AA_o_bits;
  assign AsyncQueue_3_io_deq_clock = io_clk_ARM;
  assign AsyncQueue_3_io_deq_ready = io_ARM_Flag_AA_o_ready;
  assign AsyncQueue_4_io_enq_clock = io_clk_PDA;
  assign AsyncQueue_4_io_enq_valid = ble_packetdisassembler_io_DMA_Flag_CRC_o_valid;
  assign AsyncQueue_4_io_enq_bits = ble_packetdisassembler_io_DMA_Flag_CRC_o_bits;
  assign AsyncQueue_4_io_deq_clock = io_clk_ARM;
  assign AsyncQueue_4_io_deq_ready = io_ARM_Flag_CRC_o_ready;
endmodule
